module ARR_CONTROLLER(
    input clk,
    input rstn,
    input config_dat_in,
    input config_num_in,

)