* SPICE NETLIST
***************************************

.SUBCKT esdscr A K PD SX
.ENDS
***************************************
.SUBCKT subc SUBCON SUB
.ENDS
***************************************
.SUBCKT sblkndres D S G
.ENDS
***************************************
.SUBCKT ncap G S B D
.ENDS
***************************************
.SUBCKT dgncap G S B D
.ENDS
***************************************
.SUBCKT diffhavar ANODE1 ANODE2 CATHODE BULK
.ENDS
***************************************
.SUBCKT diffncap GA GB NW SX
.ENDS
***************************************
.SUBCKT esdnsh_base d g s b
.ENDS
***************************************
.SUBCKT esdpsh_base d g s b
.ENDS
***************************************
.SUBCKT bondpad in gp sub
.ENDS
***************************************
.SUBCKT devicepad pad
.ENDS
***************************************
.SUBCKT efuse IN OUT
.ENDS
***************************************
.SUBCKT indp out in bulk
.ENDS
***************************************
.SUBCKT ind out in bulk
.ENDS
***************************************
.SUBCKT inds out in bulk
.ENDS
***************************************
.SUBCKT symindp outpr outse ct BULK
.ENDS
***************************************
.SUBCKT symind outpr outse ct BULK
.ENDS
***************************************
.SUBCKT rfline in out bulk
.ENDS
***************************************
.SUBCKT singlewire VA VB VSHIELD
.ENDS
***************************************
.SUBCKT coupledwires VA1 VA2 VB1 VB2 VSHIELD
.ENDS
***************************************
.SUBCKT singlecpw va vb vshield
.ENDS
***************************************
.SUBCKT coupledcpw va1 va2 vb1 vb2 vshield
.ENDS
***************************************
.SUBCKT corrPoint cp
.ENDS
***************************************
.SUBCKT FILL1TS
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT FILL2TS
** N=6 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_1
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT INVX1TS
** N=14 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VSS VDD A Y
.ENDS
***************************************
.SUBCKT NOR2X1TS
** N=20 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B VDD A Y VSS
.ENDS
***************************************
.SUBCKT FILL4TS
** N=10 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_2
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT INVX2TS
** N=14 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A VSS VDD Y
.ENDS
***************************************
.SUBCKT OR2X1TS
** N=25 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VSS A B VDD Y
.ENDS
***************************************
.SUBCKT NAND2BX2TS
** N=31 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: AN B VDD Y VSS
.ENDS
***************************************
.SUBCKT NOR2BX2TS
** N=34 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: AN B Y VSS VDD
.ENDS
***************************************
.SUBCKT FILL8TS
** N=18 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT CLKAND2X2TS
** N=23 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A B VSS VDD Y
.ENDS
***************************************
.SUBCKT NOR2X2TS
** N=26 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A B Y VSS VDD
.ENDS
***************************************
.SUBCKT AOI21X4TS
** N=48 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A0 A1 VDD B0 VSS Y
.ENDS
***************************************
.SUBCKT AOI21X2TS
** N=43 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A1 VDD A0 B0 VSS Y
.ENDS
***************************************
.SUBCKT OR2X2TS
** N=26 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A B VSS VDD Y
.ENDS
***************************************
.SUBCKT NAND2X1TS
** N=19 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B VSS Y A VDD
.ENDS
***************************************
.SUBCKT NOR2BX1TS
** N=25 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: AN B VDD Y VSS
.ENDS
***************************************
.SUBCKT XNOR2X4TS
** N=64 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B A Y VSS VDD
.ENDS
***************************************
.SUBCKT XOR2X4TS
** N=74 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B A Y VSS VDD
.ENDS
***************************************
.SUBCKT NAND2X2TS
** N=26 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VSS A B Y VDD
.ENDS
***************************************
.SUBCKT ICV_3
** N=8 EP=0 IP=10 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT OAI2BB1X2TS
** N=37 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A1N A0N Y B0 VDD VSS
.ENDS
***************************************
.SUBCKT AND2X2TS
** N=26 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A B VDD VSS Y
.ENDS
***************************************
.SUBCKT OAI21XLTS
** N=23 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A1 VSS A0 B0 VDD Y
.ENDS
***************************************
.SUBCKT DFFRHQX2TS
** N=94 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: CK D RN VDD VSS Q
.ENDS
***************************************
.SUBCKT FILL16TS
** N=36 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT AO22XLTS
** N=35 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B1 B0 A0 A1 VDD VSS Y
.ENDS
***************************************
.SUBCKT DFFRXLTS
** N=85 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: D CK RN QN VDD VSS Q
.ENDS
***************************************
.SUBCKT OAI21X1TS
** N=24 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A1 VSS A0 B0 VDD Y
.ENDS
***************************************
.SUBCKT FILL32TS
** N=74 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT CLKINVX2TS
** N=14 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A VSS VDD Y
.ENDS
***************************************
.SUBCKT INVX6TS
** N=24 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A VSS Y VDD
.ENDS
***************************************
.SUBCKT ICV_4
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT OAI21X2TS
** N=45 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A0 A1 VSS B0 Y VDD
.ENDS
***************************************
.SUBCKT NOR2X4TS
** N=36 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B VDD A VSS Y
.ENDS
***************************************
.SUBCKT NOR2XLTS
** N=20 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B VDD A Y VSS
.ENDS
***************************************
.SUBCKT AOI21X1TS
** N=24 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A1 A0 VDD B0 VSS Y
.ENDS
***************************************
.SUBCKT BUFX4TS
** N=27 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A Y VSS VDD
.ENDS
***************************************
.SUBCKT CLKBUFX2TS
** N=18 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A VSS VDD Y
.ENDS
***************************************
.SUBCKT BUFX3TS
** N=21 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A Y VSS VDD
.ENDS
***************************************
.SUBCKT ICV_5
** N=6 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT DFFRHQX4TS
** N=113 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: CK D RN Q VSS VDD
.ENDS
***************************************
.SUBCKT ICV_6
** N=8 EP=0 IP=10 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_7
** N=43 EP=0 IP=46 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT NAND2BX1TS
** N=22 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: AN B VSS Y VDD
.ENDS
***************************************
.SUBCKT INVX4TS
** N=19 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A Y VSS VDD
.ENDS
***************************************
.SUBCKT OAI21X4TS
** N=47 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A1 VSS A0 B0 Y VDD
.ENDS
***************************************
.SUBCKT INVX8TS
** N=28 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A Y VDD VSS
.ENDS
***************************************
.SUBCKT XNOR2X2TS
** N=50 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B A VSS VDD Y
.ENDS
***************************************
.SUBCKT NAND2X4TS
** N=30 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B VSS A Y VDD
.ENDS
***************************************
.SUBCKT NAND2X6TS
** N=42 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A B Y VDD VSS
.ENDS
***************************************
.SUBCKT NOR2BX4TS
** N=38 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: AN B VDD VSS Y
.ENDS
***************************************
.SUBCKT OR2X4TS
** N=32 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A B Y VDD VSS
.ENDS
***************************************
.SUBCKT INVX3TS
** N=20 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A Y VDD VSS
.ENDS
***************************************
.SUBCKT CMPR32X2TS
** N=81 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B A C CO VSS VDD S
.ENDS
***************************************
.SUBCKT OAI22X2TS
** N=50 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B0 VSS B1 A0 Y A1 VDD
.ENDS
***************************************
.SUBCKT DFFRX1TS
** N=85 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: D CK RN QN VDD VSS Q
.ENDS
***************************************
.SUBCKT ADDFHX2TS
** N=111 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A B CI CO VSS VDD S
.ENDS
***************************************
.SUBCKT OA21X4TS
** N=45 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A1 A0 B0 VDD Y VSS
.ENDS
***************************************
.SUBCKT OAI22X1TS
** N=32 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B1 VSS B0 A0 A1 VDD Y
.ENDS
***************************************
.SUBCKT OAI22X4TS
** N=53 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B0 B1 VSS A1 VDD A0 Y
.ENDS
***************************************
.SUBCKT AO21X2TS
** N=34 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A1 A0 B0 VSS VDD Y
.ENDS
***************************************
.SUBCKT CLKINVX4TS
** N=21 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A Y VSS VDD
.ENDS
***************************************
.SUBCKT ADDFHX4TS
** N=170 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A B CI CO S VSS VDD
.ENDS
***************************************
.SUBCKT XNOR2X1TS
** N=31 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B A Y VDD VSS
.ENDS
***************************************
.SUBCKT BUFX8TS
** N=39 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A Y VSS VDD
.ENDS
***************************************
.SUBCKT BUFX6TS
** N=36 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A VDD VSS Y
.ENDS
***************************************
.SUBCKT CLKINVX6TS
** N=27 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A VSS VDD Y
.ENDS
***************************************
.SUBCKT CLKINVX1TS
** N=13 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A VSS VDD Y
.ENDS
***************************************
.SUBCKT DFFRX2TS
** N=89 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: D CK RN VSS VDD Q QN
.ENDS
***************************************
.SUBCKT OAI2BB1X4TS
** N=40 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A1N A0N B0 VSS VDD Y
.ENDS
***************************************
.SUBCKT XOR2X1TS
** N=30 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A B Y VDD VSS
.ENDS
***************************************
.SUBCKT XOR2XLTS
** N=30 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A B Y VSS VDD
.ENDS
***************************************
.SUBCKT NAND2BX4TS
** N=41 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: AN B VSS VDD Y
.ENDS
***************************************
.SUBCKT ADDHX2TS
** N=74 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B S A VSS VDD CO
.ENDS
***************************************
.SUBCKT NAND2BXLTS
** N=23 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: AN B VSS Y VDD
.ENDS
***************************************
.SUBCKT CLKBUFX4TS
** N=31 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A Y VSS VDD
.ENDS
***************************************
.SUBCKT BUFX2TS
** N=22 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A Y VSS VDD
.ENDS
***************************************
.SUBCKT PE data_in[3] VSS data_in[0] VDD data_in[1] data_in[5] data_in[6] data_in[4] data_in[2] data_in[7] clk rst_n weight_out[0] weight_in[0] weight_in[1] weight_in[2] weight_in[3] weight_in[4] weight_in[5] weight_in[6]
+ weight_in[7] fire_in result[1] result[2] result[5] result[4] result[7] result[6] result[3] result[10] result[9] result[8] result[12] result[11] result[13] result[14] result[17] result[19] result[24] result[23]
+ result[21] result[25] result[20] result[27] result[26] result[28] result[29] result[30] result[31] data_out[0] data_out[1] data_out[2] data_out[3] data_out[4] data_out[5] data_out[6] data_out[7] weight_out[1] weight_out[2] weight_out[3]
+ weight_out[4] weight_out[5] weight_out[6] weight_out[7] fire_out result[0] result[15] result[16] result[18] result[22]
** N=4526 EP=70 IP=7193 FDC=10040
M0 946 870 872 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.4e-14 as=1.308e-13 pd=4.4e-07 ps=1.52e-06 nrd=0.416667 nrs=2.27083 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=8860 $Y=75510 $D=28
M1 947 37 946 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.4e-14 as=2.4e-14 pd=4.4e-07 ps=4.4e-07 nrd=0.416667 nrs=0.416667 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=9180 $Y=75510 $D=28
M2 VSS 32 947 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.60062e-13 as=2.4e-14 pd=1.41231e-06 ps=4.4e-07 nrd=2.77885 nrs=0.416667 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=9500 $Y=75510 $D=28
M3 VSS clk 870 VSS lpnfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26962e-13 as=1.216e-13 pd=1.23289e-06 ps=1.4e-06 nrd=0.87924 nrs=0.842105 sa=3.2e-07 sb=6.63684e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=10480 $Y=75660 $D=28
M4 VSS data_in[2] 871 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.36459e-14 as=9.6e-14 pd=5.87869e-07 ps=1.28e-06 nrd=1.52161 nrs=1.98347 sa=3.6e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=8.4e-15 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=10520 $Y=32520 $D=28
M5 874 870 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=8.01867e-14 pd=1.28e-06 ps=7.78667e-07 nrd=1.69444 nrs=1.39213 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=1.32e-14 panw8=0 panw9=0 panw10=0 $X=10990 $Y=75660 $D=28
M6 141 871 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.41023e-13 pd=2.08e-06 ps=1.92393e-06 nrd=0.444444 nrs=0.464936 sa=5.31111e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=11080 $Y=32290 $D=28
M7 949 874 872 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.46e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=12010 $Y=75590 $D=28
M8 950 873 949 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=1.14e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=12330 $Y=75590 $D=28
M9 VSS 32 950 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.8e-14 as=2e-14 pd=9.77778e-07 ps=4e-07 nrd=2.2 nrs=0.5 sa=1e-06 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=12650 $Y=75590 $D=28
M10 873 872 VSS VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.168e-13 as=1.496e-13 pd=1.08e-06 ps=1.66222e-06 nrd=1.01038 nrs=1.29412 sa=9.65882e-07 sb=4.25882e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=13110 $Y=75590 $D=28
M11 875 874 873 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48844e-13 as=1.168e-13 pd=1.42296e-06 ps=1.08e-06 nrd=1.28758 nrs=1.01038 sa=4.14118e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.2e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=13670 $Y=75890 $D=28
M12 952 870 875 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.75556e-14 pd=4e-07 ps=8.37037e-07 nrd=0.5 nrs=2.18889 sa=3.6e-07 sb=1.46e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=14230 $Y=75570 $D=28
M13 VSS 878 952 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.37333e-14 as=2e-14 pd=4.02222e-07 ps=4e-07 nrd=1.34333 nrs=0.5 sa=6.8e-07 sb=1.14e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=14550 $Y=75570 $D=28
M14 953 32 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.2e-14 as=2.47173e-13 pd=1.12e-06 ps=1.85022e-06 nrd=0.108696 nrs=0.292029 sa=5.64565e-07 sb=6.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=15030 $Y=75490 $D=28
M15 878 875 953 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=9.2e-14 pd=2.52e-06 ps=1.12e-06 nrd=0.369565 nrs=0.108696 sa=8.84565e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=15350 $Y=75490 $D=28
M16 VSS 878 876 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.06635e-13 as=1.408e-13 pd=8.54118e-07 ps=1.52e-06 nrd=0.550802 nrs=0.727273 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-15 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=16310 $Y=75970 $D=28
M17 877 876 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.22965e-13 pd=1.28e-06 ps=1.78588e-06 nrd=0.195652 nrs=0.263427 sa=5.68696e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=16830 $Y=75490 $D=28
M18 VSS 876 877 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.0487e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=17310 $Y=75490 $D=28
M19 239 878 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.5287e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=17790 $Y=75490 $D=28
M20 VSS 878 239 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=1.87478e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=18270 $Y=75490 $D=28
M21 VSS clk 879 VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.15242e-13 as=1.064e-13 pd=1.04632e-06 ps=1.32e-06 nrd=1.46992 nrs=1.35714 sa=3.6e-07 sb=7.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.28e-14 panw8=0 panw9=0 panw10=0 $X=20160 $Y=18100 $D=28
M22 882 clk VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=8.23158e-14 pd=1.28e-06 ps=7.47368e-07 nrd=2.36 nrs=2.05789 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=1.32e-14 panw8=0 panw9=0 panw10=0 $X=20720 $Y=18100 $D=28
M23 880 95 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=1.04667e-13 pd=1.28e-06 ps=1e-06 nrd=2.36 nrs=2.61667 sa=3.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.2e-15 panw8=2.28e-14 panw9=0 panw10=0 $X=21760 $Y=18240 $D=28
M24 VSS 879 884 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.17059e-14 as=1.08e-13 pd=1.06471e-06 ps=1.32e-06 nrd=1.01895 nrs=1.2 sa=3.6e-07 sb=1.595e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.2e-15 panw8=0 panw9=0 panw10=0 $X=22800 $Y=17760 $D=28
M25 956 882 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.4e-14 as=1.34502e-13 pd=6.4e-07 ps=1.56157e-06 nrd=0.227273 nrs=0.694742 sa=6.55909e-07 sb=1.25409e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=23290 $Y=17760 $D=28
M26 881 880 956 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.14812e-13 as=4.4e-14 pd=1.2375e-06 ps=6.4e-07 nrd=0.59304 nrs=0.227273 sa=9.75909e-07 sb=1.07955e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=23610 $Y=17760 $D=28
M27 958 884 881 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.21875e-14 pd=4e-07 ps=5.625e-07 nrd=0.5 nrs=1.30469 sa=1.5975e-06 sb=1.94e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=24190 $Y=17910 $D=28
M28 VSS 883 958 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.3434e-14 as=2e-14 pd=6.07547e-07 ps=4e-07 nrd=1.33585 nrs=0.5 sa=1.865e-06 sb=1.78e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=24510 $Y=17910 $D=28
M29 959 68 VSS VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.67e-14 as=1.54958e-13 pd=8.1e-07 ps=1.76189e-06 nrd=0.198276 nrs=0.460638 sa=8.38276e-07 sb=1.36241e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=24950 $Y=17910 $D=28
M30 883 881 959 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29132e-13 as=6.67e-14 pd=1.12717e-06 ps=8.1e-07 nrd=0.383865 nrs=0.198276 sa=1.07621e-06 sb=1.1331e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=25300 $Y=17910 $D=28
M31 887 884 883 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.11247e-13 as=1.06868e-13 pd=1.24235e-06 ps=9.3283e-07 nrd=0.482843 nrs=0.463836 sa=1.51e-06 sb=8.03333e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=25870 $Y=17910 $D=28
M32 960 882 887 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=4.63529e-14 pd=4e-07 ps=5.17647e-07 nrd=0.5 nrs=1.15882 sa=1.84e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=26390 $Y=18010 $D=28
M33 961 68 960 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=2e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=26710 $Y=18010 $D=28
M34 VSS 886 961 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33167e-13 as=2e-14 pd=1.20833e-06 ps=4e-07 nrd=3.32917 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=27030 $Y=18010 $D=28
M35 VSS 887 886 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.91064e-14 as=9.44e-14 pd=6.93617e-07 ps=1.28e-06 nrd=1.72766 nrs=2.36 sa=3.6e-07 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=28630 $Y=17890 $D=28
M36 100 887 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.58945e-13 pd=1.56e-06 ps=1.59532e-06 nrd=0.695652 nrs=0.751156 sa=4.83478e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=29070 $Y=17890 $D=28
M37 963 888 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.2e-14 as=2.944e-13 pd=1.12e-06 ps=2.48e-06 nrd=0.108696 nrs=0.347826 sa=3.2e-07 sb=1.80783e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=30490 $Y=69990 $D=28
M38 889 105 963 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=9.2e-14 pd=1.28e-06 ps=1.12e-06 nrd=0.195652 nrs=0.108696 sa=6.4e-07 sb=1.71739e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=30810 $Y=69990 $D=28
M39 964 105 889 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.2e-14 as=1.656e-13 pd=1.12e-06 ps=1.28e-06 nrd=0.108696 nrs=0.195652 sa=1.12e-06 sb=1.58174e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=31290 $Y=69990 $D=28
M40 VSS 888 964 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.45489e-13 as=9.2e-14 pd=1.72354e-06 ps=1.12e-06 nrd=0.290039 nrs=0.108696 sa=1.44e-06 sb=1.4913e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=31610 $Y=69990 $D=28
M41 402 889 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20972e-13 as=1.76111e-13 pd=1.06937e-06 ps=1.23646e-06 nrd=0.277714 nrs=0.404296 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=32290 $Y=70250 $D=28
M42 VSS 889 402 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.68628e-13 pd=1.28e-06 ps=1.49063e-06 nrd=0.195652 nrs=0.199229 sa=1.4913e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=32770 $Y=69990 $D=28
M43 402 889 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.62696e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=33250 $Y=69990 $D=28
M44 VSS 889 402 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=1.76261e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=33730 $Y=69990 $D=28
M45 965 890 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=2.45464e-13 pd=8.6e-07 ps=1.99404e-06 nrd=0.151515 nrs=0.563507 sa=3.6e-07 sb=1.79121e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.08e-14 panw10=0 $X=36480 $Y=68420 $D=28
M46 966 807 965 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=6.6e-14 pd=8.6e-07 ps=8.6e-07 nrd=0.151515 nrs=0.151515 sa=6.8e-07 sb=1.55152e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.08e-14 panw10=0 $X=36800 $Y=68420 $D=28
M47 190 161 966 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=6.6e-14 pd=1.17e-06 ps=8.6e-07 nrd=0.305785 nrs=0.151515 sa=1e-06 sb=1.23152e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.08e-14 panw10=0 $X=37120 $Y=68420 $D=28
M48 967 161 190 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=1.332e-13 pd=8.6e-07 ps=1.17e-06 nrd=0.151515 nrs=0.305785 sa=1.24394e-06 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=37620 $Y=68290 $D=28
M49 968 807 967 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=6.6e-14 pd=8.6e-07 ps=8.6e-07 nrd=0.151515 nrs=0.151515 sa=1.56394e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=37940 $Y=68290 $D=28
M50 VSS 890 968 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.112e-13 as=6.6e-14 pd=1.96e-06 ps=8.6e-07 nrd=0.484848 nrs=0.151515 sa=1.77152e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=38260 $Y=68290 $D=28
M51 969 147 891 VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=8.96e-14 pd=4.8e-07 ps=1.2e-06 nrd=0.357143 nrs=1.14286 sa=3.2e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=38960 $Y=17950 $D=28
M52 VSS 143 969 VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.33655e-14 as=2.8e-14 pd=7.57931e-07 ps=4.8e-07 nrd=1.19089 nrs=0.357143 sa=6.4e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=39280 $Y=17950 $D=28
M53 970 154 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.00069e-13 pd=8e-07 ps=1.62414e-06 nrd=0.166667 nrs=0.555747 sa=7.52e-07 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=39840 $Y=17950 $D=28
M54 892 153 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=40010 $Y=75490 $D=28
M55 125 891 970 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=1.072e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=40160 $Y=17950 $D=28
M56 VSS 153 892 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=40490 $Y=75490 $D=28
M57 135 892 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.28e-06 sb=1.9113e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=40970 $Y=75490 $D=28
M58 VSS 892 135 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.76e-06 sb=1.73391e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=41450 $Y=75490 $D=28
M59 135 892 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=2e-06 sb=1.46196e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=41930 $Y=75490 $D=28
M60 VSS 892 135 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.09024e-13 as=1.656e-13 pd=1.6192e-06 ps=1.28e-06 nrd=0.246957 nrs=0.195652 sa=2e-06 sb=9.81957e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=42410 $Y=75490 $D=28
M61 135 892 VSS VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.044e-13 as=1.31776e-13 pd=9.4e-07 ps=1.0208e-06 nrd=0.310345 nrs=0.391724 sa=2e-06 sb=8.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=9.6e-15 panw9=0 panw10=0 $X=42930 $Y=75490 $D=28
M62 VSS 892 135 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.146e-13 as=1.044e-13 pd=1.9e-06 ps=9.4e-07 nrd=0.637931 nrs=0.310345 sa=2e-06 sb=3.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=9.6e-15 panw9=0 panw10=0 $X=43410 $Y=75490 $D=28
M63 VSS 897 896 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.55477e-13 as=2.944e-13 pd=1.92256e-06 ps=2.48e-06 nrd=0.301839 nrs=0.347826 sa=3.2e-07 sb=5.6087e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=60040 $Y=25090 $D=28
M64 895 227 VSS VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=9.99692e-14 pd=1.36e-06 ps=7.52308e-07 nrd=0.888889 nrs=0.771368 sa=8.8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=60600 $Y=25210 $D=28
M65 244 895 896 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.764e-13 pd=1.28e-06 ps=2.8e-06 nrd=0.195652 nrs=0.32656 sa=3.00435e-07 sb=1.6638e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=61780 $Y=25090 $D=28
M66 897 227 244 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.68875e-13 as=1.656e-13 pd=1.33062e-06 ps=1.28e-06 nrd=0.199521 nrs=0.195652 sa=7.80435e-07 sb=1.27511e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=62260 $Y=25090 $D=28
M67 VSS 264 897 VSS lpnfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99561e-13 as=1.56025e-13 pd=1.615e-06 ps=1.22938e-06 nrd=0.276209 nrs=0.215952 sa=1.26871e-06 sb=8.77882e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=62740 $Y=25160 $D=28
M68 901 195 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.7759e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.587076 sa=2.4e-07 sb=1.94e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=63170 $Y=46690 $D=28
M69 897 264 VSS VSS lpnfet w=4.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.196e-13 as=1.00954e-13 pd=1.5e-06 ps=8.17e-07 nrd=0.646836 nrs=0.545995 sa=1.72e-06 sb=2.7814e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=63300 $Y=25160 $D=28
M70 971 264 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.2e-14 as=5.63467e-14 pd=5.9e-07 ps=4.56e-07 nrd=0.729167 nrs=0.978241 sa=2e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=2.64e-14 panw10=0 $X=63300 $Y=25770 $D=28
M71 VSS 195 901 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=7.2e-07 sb=1.636e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=63650 $Y=46690 $D=28
M72 898 227 971 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=4.2e-14 pd=1.28e-06 ps=5.9e-07 nrd=1.69444 nrs=0.729167 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=2.64e-14 panw10=0 $X=63770 $Y=25770 $D=28
M73 900 901 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.155e-13 as=1.24348e-13 pd=9.7e-07 ps=1.29928e-06 nrd=0.381818 nrs=0.411067 sa=1.16e-06 sb=1.196e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=64090 $Y=46690 $D=28
M74 VSS 898 205 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7107e-13 as=1.472e-13 pd=1.92703e-06 ps=1.56e-06 nrd=0.808461 nrs=0.695652 sa=3.2e-07 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=64350 $Y=25090 $D=28
M75 VSS 901 900 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28174e-13 as=1.155e-13 pd=1.19565e-06 ps=9.7e-07 nrd=0.423715 nrs=0.381818 sa=1.7e-06 sb=6.56e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=64630 $Y=46690 $D=28
M76 899 187 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02539e-13 pd=1.52e-06 ps=9.56522e-07 nrd=0.727273 nrs=0.529644 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=65070 $Y=46690 $D=28
M77 900 899 245 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.544e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.510413 sa=2.80727e-07 sb=1.57455e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=8.4e-15 panw9=0 panw10=0 $X=66030 $Y=46710 $D=28
M78 903 906 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.22478e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=66210 $Y=62790 $D=28
M79 245 899 900 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07578e-13 as=9.9e-14 pd=1.00917e-06 ps=9.1e-07 nrd=0.35563 nrs=0.327273 sa=7.60727e-07 sb=1.09455e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=8.4e-15 panw9=0 panw10=0 $X=66510 $Y=46710 $D=28
M80 VSS 906 903 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.22525e-13 as=1.656e-13 pd=1.56208e-06 ps=1.28e-06 nrd=0.262908 nrs=0.195652 sa=8e-07 sb=7.44783e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=66690 $Y=62790 $D=28
M81 901 187 245 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.72e-14 as=1.05622e-13 pd=9e-07 ps=9.90826e-07 nrd=0.333333 nrs=0.362215 sa=1.07333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=66990 $Y=46810 $D=28
M82 902 266 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.1e-13 as=1.7415e-13 pd=2.08e-06 ps=1.2225e-06 nrd=0.405093 nrs=0.335937 sa=1.36e-06 sb=2.91667e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=67250 $Y=62990 $D=28
M83 245 187 901 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=9.72e-14 pd=1.72e-06 ps=9e-07 nrd=0.592593 nrs=0.333333 sa=1.55333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=67470 $Y=46810 $D=28
M84 903 902 250 VSS lpnfet w=8.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.494e-13 as=2.656e-13 pd=1.19e-06 ps=2.3e-06 nrd=0.216867 nrs=0.385542 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=68350 $Y=62790 $D=28
M85 250 902 903 VSS lpnfet w=8.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.49885e-13 as=1.494e-13 pd=1.20374e-06 ps=1.19e-06 nrd=0.217572 nrs=0.216867 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=68830 $Y=62790 $D=28
M86 906 266 250 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.584e-13 as=1.58915e-13 pd=1.24e-06 ps=1.27626e-06 nrd=0.204545 nrs=0.20521 sa=1.21864e-06 sb=8e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=69310 $Y=62790 $D=28
M87 250 266 906 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=1.584e-13 pd=2.4e-06 ps=1.24e-06 nrd=0.363636 nrs=0.204545 sa=1.69864e-06 sb=3.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=69790 $Y=62790 $D=28
M88 972 266 905 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.8e-14 as=1.536e-13 pd=6.8e-07 ps=1.6e-06 nrd=0.208333 nrs=0.666667 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=70730 $Y=63200 $D=28
M89 VSS 260 972 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8827e-14 as=4.8e-14 pd=9.42331e-07 ps=6.8e-07 nrd=0.428937 nrs=0.208333 sa=6.4e-07 sb=1.8e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=71050 $Y=63200 $D=28
M90 906 260 VSS VSS lpnfet w=8.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.566e-13 as=1.79124e-13 pd=1.23e-06 ps=1.70798e-06 nrd=0.206897 nrs=0.236655 sa=7.11724e-07 sb=1.34207e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=71490 $Y=62810 $D=28
M91 VSS 260 906 VSS lpnfet w=8.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.01805e-13 as=1.566e-13 pd=1.39899e-06 ps=1.23e-06 nrd=0.26662 nrs=0.206897 sa=1.19172e-06 sb=8.62069e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=71970 $Y=62810 $D=28
M92 906 260 VSS VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.94846e-13 pd=2.32e-06 ps=1.35075e-06 nrd=0.380952 nrs=0.276143 sa=1.69571e-06 sb=3.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=72530 $Y=62840 $D=28
M93 276 905 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.944e-13 pd=2.48e-06 ps=2.48e-06 nrd=0.347826 nrs=0.347826 sa=3.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=73470 $Y=62790 $D=28
M94 353 323 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=3.78986e-13 pd=1.22e-06 ps=1.84705e-06 nrd=0.209302 nrs=0.512421 sa=7.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=85760 $Y=75550 $D=28
M95 974 301 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.4e-14 as=1.056e-13 pd=4.4e-07 ps=1.34e-06 nrd=0.416667 nrs=1.83333 sa=3.7e-07 sb=1.555e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=86060 $Y=39640 $D=28
M96 VSS 342 353 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9522e-13 as=1.548e-13 pd=1.3502e-06 ps=1.22e-06 nrd=0.263953 nrs=0.209302 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=86240 $Y=75550 $D=28
M97 908 232 974 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.41818e-14 as=2.4e-14 pd=8.72727e-07 ps=4.4e-07 nrd=1.28788 nrs=0.416667 sa=6.9e-07 sb=1.235e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=86380 $Y=39640 $D=28
M98 353 342 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=1.9522e-13 pd=1.22e-06 ps=1.3502e-06 nrd=0.209302 nrs=0.263953 sa=1.8e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=86800 $Y=75550 $D=28
M99 VSS 314 908 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.59574e-14 as=6.18182e-14 pd=6.97872e-07 ps=7.27273e-07 nrd=1.89894 nrs=1.54545 sa=1.25e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=6e-15 panw8=0 panw9=0 panw10=0 $X=86940 $Y=39640 $D=28
M100 VSS 323 353 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9522e-13 as=1.548e-13 pd=1.3502e-06 ps=1.22e-06 nrd=0.263953 nrs=0.209302 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=87280 $Y=75550 $D=28
M101 413 908 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.74702e-13 pd=1.56e-06 ps=1.60511e-06 nrd=0.695652 nrs=0.825624 sa=9.60435e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=87470 $Y=39490 $D=28
M102 353 323 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=1.9522e-13 pd=1.22e-06 ps=1.3502e-06 nrd=0.209302 nrs=0.263953 sa=2e-06 sb=1.88e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=87840 $Y=75550 $D=28
M103 VSS 342 353 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9522e-13 as=1.548e-13 pd=1.3502e-06 ps=1.22e-06 nrd=0.263953 nrs=0.209302 sa=2e-06 sb=1.4e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=88320 $Y=75550 $D=28
M104 353 342 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=1.9522e-13 pd=1.22e-06 ps=1.3502e-06 nrd=0.209302 nrs=0.263953 sa=2e-06 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=88880 $Y=75550 $D=28
M105 VSS 323 353 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.90589e-13 as=1.548e-13 pd=2.24807e-06 ps=1.22e-06 nrd=0.392901 nrs=0.209302 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=89360 $Y=75550 $D=28
M106 979 375 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.8e-14 as=2.816e-13 pd=1.08e-06 ps=2.4e-06 nrd=0.113636 nrs=0.363636 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=102820 $Y=61120 $D=28
M107 980 379 979 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.8e-14 as=8.8e-14 pd=1.08e-06 ps=1.08e-06 nrd=0.113636 nrs=0.113636 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=103140 $Y=61120 $D=28
M108 382 391 980 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.584e-13 as=8.8e-14 pd=1.24e-06 ps=1.08e-06 nrd=0.204545 nrs=0.113636 sa=9.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=103460 $Y=61120 $D=28
M109 981 391 382 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.8e-14 as=1.584e-13 pd=1.08e-06 ps=1.24e-06 nrd=0.113636 nrs=0.204545 sa=1.44e-06 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=103940 $Y=61120 $D=28
M110 982 379 981 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.8e-14 as=8.8e-14 pd=1.08e-06 ps=1.08e-06 nrd=0.113636 nrs=0.113636 sa=1.76e-06 sb=1.89955e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=104260 $Y=61120 $D=28
M111 VSS 375 982 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00847e-13 as=8.8e-14 pd=1.38039e-06 ps=1.08e-06 nrd=0.259358 nrs=0.113636 sa=2e-06 sb=1.57955e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=104580 $Y=61120 $D=28
M112 983 375 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.8e-14 as=2.00847e-13 pd=1.08e-06 ps=1.38039e-06 nrd=0.113636 nrs=0.259358 sa=2e-06 sb=1.01955e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=105140 $Y=61120 $D=28
M113 984 379 983 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.8e-14 as=8.8e-14 pd=1.08e-06 ps=1.08e-06 nrd=0.113636 nrs=0.113636 sa=2e-06 sb=6.99545e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=105460 $Y=61120 $D=28
M114 382 391 984 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.34e-13 as=8.8e-14 pd=2.56e-06 ps=1.08e-06 nrd=0.431302 nrs=0.113636 sa=2e-06 sb=3.79545e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=105780 $Y=61120 $D=28
M115 417 401 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-15 $X=106020 $Y=69990 $D=28
M116 VSS 392 417 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=6e-15 $X=106500 $Y=69990 $D=28
M117 417 392 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=6e-15 $X=106980 $Y=69990 $D=28
M118 VSS 401 417 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.76e-06 sb=1.72e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=6e-15 $X=107460 $Y=69990 $D=28
M119 417 401 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=2e-06 sb=1.24e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=6e-15 $X=107940 $Y=69990 $D=28
M120 VSS 392 417 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.15112e-13 as=1.656e-13 pd=1.97143e-06 ps=1.28e-06 nrd=0.490444 nrs=0.195652 sa=2e-06 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=108420 $Y=69990 $D=28
M121 911 448 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=119240 $Y=55960 $D=28
M122 VSS 433 911 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=119720 $Y=55960 $D=28
M123 911 433 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=120200 $Y=55960 $D=28
M124 VSS 448 911 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12844e-13 as=9.9e-14 pd=9.57823e-07 ps=9.1e-07 nrd=0.373036 nrs=0.327273 sa=1.76e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=120680 $Y=55960 $D=28
M125 443 911 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.88756e-13 pd=1.28e-06 ps=1.60218e-06 nrd=0.195652 nrs=0.223011 sa=1.30826e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=121160 $Y=55590 $D=28
M126 VSS 911 443 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.5013e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=121640 $Y=55590 $D=28
M127 443 911 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=1.69435e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=122120 $Y=55590 $D=28
M128 545 523 VSS VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.46e-14 as=1.61e-13 pd=8.3e-07 ps=1.64e-06 nrd=0.382979 nrs=0.728837 sa=3.42553e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=134910 $Y=54270 $D=28
M129 VSS 523 545 VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.46e-14 as=8.46e-14 pd=8.3e-07 ps=8.3e-07 nrd=0.382979 nrs=0.382979 sa=8.22553e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=135390 $Y=54270 $D=28
M130 545 523 VSS VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.46e-14 as=8.46e-14 pd=8.3e-07 ps=8.3e-07 nrd=0.382979 nrs=0.382979 sa=1.30255e-06 sb=1.88e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=135870 $Y=54270 $D=28
M131 VSS 523 545 VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16344e-13 as=8.46e-14 pd=9.63115e-07 ps=8.3e-07 nrd=0.526683 nrs=0.382979 sa=1.78255e-06 sb=1.4e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=136350 $Y=54270 $D=28
M132 545 523 VSS VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.46e-14 as=1.16344e-13 pd=8.3e-07 ps=9.63115e-07 nrd=0.382979 nrs=0.526683 sa=2e-06 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=136910 $Y=54270 $D=28
M133 VSS 523 545 VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.65691e-13 as=8.46e-14 pd=1.4664e-06 ps=8.3e-07 nrd=0.750071 nrs=0.382979 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=137390 $Y=54270 $D=28
M134 991 608 915 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.4e-14 as=2.236e-13 pd=4.4e-07 ps=2.18e-06 nrd=0.416667 nrs=3.88194 sa=3.6e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=139650 $Y=63350 $D=28
M135 VSS 556 991 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.11806e-13 as=2.4e-14 pd=9.05143e-07 ps=4.4e-07 nrd=1.94107 nrs=0.416667 sa=6.8e-07 sb=9.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=139970 $Y=63350 $D=28
M136 548 915 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=2.14294e-13 pd=1.56e-06 ps=1.73486e-06 nrd=0.695652 nrs=1.01273 sa=9.17391e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=140640 $Y=63250 $D=28
M137 VSS 567 916 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.06267e-13 as=1.472e-13 pd=1.08e-06 ps=1.56e-06 nrd=0.502205 nrs=0.695652 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=141610 $Y=63240 $D=28
M138 992 553 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.4e-14 as=1.47849e-13 pd=8.4e-07 ps=1.50261e-06 nrd=0.15625 nrs=0.36096 sa=6.1375e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.8e-14 panw9=0 panw10=0 $X=142050 $Y=63060 $D=28
M139 993 854 992 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.4e-14 as=6.4e-14 pd=8.4e-07 ps=8.4e-07 nrd=0.15625 nrs=0.15625 sa=9.3375e-07 sb=1.82e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.8e-14 panw9=0 panw10=0 $X=142370 $Y=63060 $D=28
M140 561 916 993 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=6.4e-14 pd=1e-06 ps=8.4e-07 nrd=0.28125 nrs=0.15625 sa=1.25375e-06 sb=1.5e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.8e-14 panw9=0 panw10=0 $X=142690 $Y=63060 $D=28
M141 994 916 561 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.4e-14 as=1.152e-13 pd=8.4e-07 ps=1e-06 nrd=0.15625 nrs=0.28125 sa=1.73375e-06 sb=1.02e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.8e-14 panw9=0 panw10=0 $X=143170 $Y=63060 $D=28
M142 995 854 994 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.4e-14 as=6.4e-14 pd=8.4e-07 ps=8.4e-07 nrd=0.15625 nrs=0.15625 sa=1.91e-06 sb=7e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.8e-14 panw9=0 panw10=0 $X=143490 $Y=63060 $D=28
M143 VSS 553 995 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.75881e-13 as=6.4e-14 pd=2.12426e-06 ps=8.4e-07 nrd=0.673537 nrs=0.15625 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.8e-14 panw9=0 panw10=0 $X=143810 $Y=63060 $D=28
M144 VSS 778 917 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.152e-13 pd=8.59701e-07 ps=1.36e-06 nrd=0.777778 nrs=0.888889 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=181440 $Y=41600 $D=28
M145 917 757 VSS VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.48e-14 as=1.008e-13 pd=7.2e-07 ps=8.59701e-07 nrd=0.5 nrs=0.777778 sa=8.8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=182000 $Y=41600 $D=28
M146 VSS 759 917 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.49846e-14 as=6.48e-14 pd=7.52308e-07 ps=7.2e-07 nrd=0.732906 nrs=0.5 sa=1.36e-06 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=182480 $Y=41600 $D=28
M147 867 917 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.42738e-13 pd=2.48e-06 ps=1.92256e-06 nrd=0.347826 nrs=0.286789 sa=9.44348e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=183040 $Y=41190 $D=28
M148 998 716 VSS VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4e-14 as=1.56e-13 pd=6e-07 ps=1.58e-06 nrd=0.25 nrs=0.975 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=183280 $Y=17940 $D=28
M149 772 765 998 VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28e-13 as=4e-14 pd=1.44e-06 ps=6e-07 nrd=0.8 nrs=0.25 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=183600 $Y=17940 $D=28
M150 137 119 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=34920 $Y=20050 $D=28
M151 270 820 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=68120 $Y=39490 $D=28
M152 821 268 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=69320 $Y=75490 $D=28
M153 387 366 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=100520 $Y=75490 $D=28
M154 471 474 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=125720 $Y=27250 $D=28
M155 465 476 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=125720 $Y=68290 $D=28
M156 478 506 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=126520 $Y=34450 $D=28
M157 484 477 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=126920 $Y=27250 $D=28
M158 489 488 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=128520 $Y=39490 $D=28
M159 486 505 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=130920 $Y=32290 $D=28
M160 547 519 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=134920 $Y=39490 $D=28
M161 531 530 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=136120 $Y=39490 $D=28
M162 914 536 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=139320 $Y=32290 $D=28
M163 550 554 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=142520 $Y=32290 $D=28
M164 529 568 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=143720 $Y=27250 $D=28
M165 565 557 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=144120 $Y=56050 $D=28
M166 572 566 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=145320 $Y=56050 $D=28
M167 603 614 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=153320 $Y=61090 $D=28
M168 630 597 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=153720 $Y=41650 $D=28
M169 601 624 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=154120 $Y=53890 $D=28
M170 639 646 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=154920 $Y=41650 $D=28
M171 619 616 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=155320 $Y=53890 $D=28
M172 635 633 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=158120 $Y=53890 $D=28
M173 642 666 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=160520 $Y=46690 $D=28
M174 648 673 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=160920 $Y=56050 $D=28
M175 670 652 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=162120 $Y=68290 $D=28
M176 640 687 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=163320 $Y=61090 $D=28
M177 675 683 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=165720 $Y=32290 $D=28
M178 698 679 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=166520 $Y=61090 $D=28
M179 862 692 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=169720 $Y=68290 $D=28
M180 759 690 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=171720 $Y=41650 $D=28
M181 720 731 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=173320 $Y=34450 $D=28
M182 709 717 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=173720 $Y=32290 $D=28
M183 677 686 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=174120 $Y=70450 $D=28
M184 757 712 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=175320 $Y=41650 $D=28
M185 750 726 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=176520 $Y=41650 $D=28
M186 728 725 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=176520 $Y=56050 $D=28
M187 730 636 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=178120 $Y=70450 $D=28
M188 748 716 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=178520 $Y=20050 $D=28
M189 765 733 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=182120 $Y=17890 $D=28
M190 707 783 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=184120 $Y=70450 $D=28
M191 773 736 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=184920 $Y=53890 $D=28
M192 918 723 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=185720 $Y=27250 $D=28
M193 776 785 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=186120 $Y=70450 $D=28
M194 786 784 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=187320 $Y=70450 $D=28
M195 422 417 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=112480 $Y=70400 $D=28
M196 VSS 431 422 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=112960 $Y=70400 $D=28
M197 438 430 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=116880 $Y=61140 $D=28
M198 VSS 437 438 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=117360 $Y=61140 $D=28
M199 458 456 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=120880 $Y=32340 $D=28
M200 VSS 471 458 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=121360 $Y=32340 $D=28
M201 472 458 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=124880 $Y=34400 $D=28
M202 VSS 489 472 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=125360 $Y=34400 $D=28
M203 488 492 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=129680 $Y=39540 $D=28
M204 VSS 497 488 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=130160 $Y=39540 $D=28
M205 516 528 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=130880 $Y=34400 $D=28
M206 VSS 519 516 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=131360 $Y=34400 $D=28
M207 510 522 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=132080 $Y=32340 $D=28
M208 VSS 509 510 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=132560 $Y=32340 $D=28
M209 528 505 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=135680 $Y=27200 $D=28
M210 VSS 529 528 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=136160 $Y=27200 $D=28
M211 539 559 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=136480 $Y=63200 $D=28
M212 VSS 608 539 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=136960 $Y=63200 $D=28
M213 549 556 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=140480 $Y=61140 $D=28
M214 VSS 608 549 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=140960 $Y=61140 $D=28
M215 581 597 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=148480 $Y=56000 $D=28
M216 VSS 588 581 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=148960 $Y=56000 $D=28
M217 673 626 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=156480 $Y=53940 $D=28
M218 VSS 624 673 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=156960 $Y=53940 $D=28
M219 666 632 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=160080 $Y=41600 $D=28
M220 VSS 639 666 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=160560 $Y=41600 $D=28
M221 686 617 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=168080 $Y=68340 $D=28
M222 VSS 657 686 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=168560 $Y=68340 $D=28
M223 703 726 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=169280 $Y=39540 $D=28
M224 VSS 675 703 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=169760 $Y=39540 $D=28
M225 685 863 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=172880 $Y=56000 $D=28
M226 VSS 695 685 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=173360 $Y=56000 $D=28
M227 710 703 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=174080 $Y=48800 $D=28
M228 VSS 713 710 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=174560 $Y=48800 $D=28
M229 745 686 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=176480 $Y=70400 $D=28
M230 VSS 730 745 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=176960 $Y=70400 $D=28
M231 737 731 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=177680 $Y=41600 $D=28
M232 VSS 712 737 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=178160 $Y=41600 $D=28
M233 783 652 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=179280 $Y=63200 $D=28
M234 VSS 744 783 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=179760 $Y=63200 $D=28
M235 788 759 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=185680 $Y=39540 $D=28
M236 VSS 778 788 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=186160 $Y=39540 $D=28
M237 769 783 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.61e-13 pd=8.2e-07 ps=1.62e-06 nrd=0.391304 nrs=0.76087 sa=3.5e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=187280 $Y=61140 $D=28
M238 VSS 785 769 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=8.28e-14 pd=2.24e-06 ps=8.2e-07 nrd=1.26276 nrs=0.391304 sa=8.3e-07 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=187760 $Y=61140 $D=28
M239 13 63 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-15 $X=14120 $Y=48390 $D=28
M240 42 52 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=16520 $Y=32290 $D=28
M241 48 43 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=17320 $Y=53890 $D=28
M242 46 133 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=17720 $Y=19590 $D=28
M243 60 58 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=20120 $Y=68290 $D=28
M244 67 81 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=24520 $Y=75490 $D=28
M245 888 885 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=29320 $Y=69990 $D=28
M246 128 117 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=34920 $Y=12390 $D=28
M247 145 893 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=41320 $Y=33990 $D=28
M248 193 181 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=48920 $Y=55590 $D=28
M249 208 815 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=56920 $Y=17890 $D=28
M250 219 237 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=58920 $Y=39490 $D=28
M251 222 230 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=62920 $Y=62790 $D=28
M252 818 215 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=64120 $Y=61090 $D=28
M253 262 249 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=68920 $Y=25090 $D=28
M254 823 272 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=70520 $Y=75490 $D=28
M255 336 284 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=78520 $Y=39490 $D=28
M256 310 339 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=82920 $Y=12390 $D=28
M257 317 363 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=85720 $Y=55590 $D=28
M258 326 339 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=91320 $Y=12390 $D=28
M259 339 345 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=91320 $Y=17890 $D=28
M260 393 376 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=103320 $Y=75490 $D=28
M261 416 380 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=107320 $Y=53890 $D=28
M262 431 473 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=113320 $Y=75490 $D=28
M263 429 417 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=115320 $Y=69990 $D=28
M264 450 427 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=119720 $Y=32290 $D=28
M265 469 458 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=123720 $Y=33990 $D=28
M266 462 844 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=125320 $Y=62790 $D=28
M267 515 509 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=127720 $Y=33990 $D=28
M268 493 456 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=131320 $Y=41190 $D=28
M269 524 497 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=131320 $Y=46690 $D=28
M270 850 479 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=134120 $Y=12390 $D=28
M271 564 850 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=140120 $Y=17890 $D=28
M272 594 523 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=144920 $Y=48390 $D=28
M273 575 586 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=145720 $Y=61090 $D=28
M274 592 586 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=149320 $Y=53890 $D=28
M275 599 607 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=152920 $Y=55590 $D=28
M276 622 617 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=156120 $Y=55590 $D=28
M277 651 655 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=163320 $Y=25090 $D=28
M278 657 576 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=163320 $Y=68290 $D=28
M279 760 658 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=164520 $Y=32290 $D=28
M280 671 703 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=165720 $Y=41190 $D=28
M281 689 860 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=169320 $Y=32290 $D=28
M282 696 695 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=174520 $Y=68290 $D=28
M283 747 734 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=179720 $Y=55590 $D=28
M284 771 867 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=184520 $Y=39490 $D=28
M285 756 918 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-14 $X=186920 $Y=26790 $D=28
M286 1727 298 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.64e-14 as=1.14542e-13 pd=8e-07 ps=1.15833e-06 nrd=1.66 nrs=2.86354 sa=3.1e-07 sb=1.35e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=74810 $Y=20150 $D=28
M287 VSS 274 1727 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.6e-14 as=6.64e-14 pd=4.94656e-07 ps=8e-07 nrd=1.15 nrs=1.66 sa=8.7e-07 sb=7.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=75370 $Y=20150 $D=28
M288 825 1727 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.058e-13 pd=1.56e-06 ps=1.13771e-06 nrd=0.695652 nrs=0.5 sa=7.35217e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=75840 $Y=19890 $D=28
M289 1729 569 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.64e-14 as=1.14542e-13 pd=8e-07 ps=1.15833e-06 nrd=1.66 nrs=2.86354 sa=3.1e-07 sb=1.35e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=144810 $Y=25250 $D=28
M290 VSS 568 1729 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.6e-14 as=6.64e-14 pd=4.94656e-07 ps=8e-07 nrd=1.15 nrs=1.66 sa=8.7e-07 sb=7.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=145370 $Y=25250 $D=28
M291 558 1729 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.058e-13 pd=1.56e-06 ps=1.13771e-06 nrd=0.695652 nrs=0.5 sa=7.35217e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=145840 $Y=25250 $D=28
M292 1731 765 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.64e-14 as=1.14542e-13 pd=8e-07 ps=1.15833e-06 nrd=1.66 nrs=2.86354 sa=3.1e-07 sb=1.35e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=186810 $Y=18050 $D=28
M293 VSS 716 1731 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.6e-14 as=6.64e-14 pd=4.94656e-07 ps=8e-07 nrd=1.15 nrs=1.66 sa=8.7e-07 sb=7.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=187370 $Y=18050 $D=28
M294 770 1731 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.058e-13 pd=1.56e-06 ps=1.13771e-06 nrd=0.695652 nrs=0.5 sa=7.35217e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=187840 $Y=18050 $D=28
M295 VSS 129 1733 VSS lpnfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02776e-13 as=1.344e-13 pd=8.56471e-07 ps=1.48e-06 nrd=0.582633 nrs=0.761905 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=55780 $Y=32290 $D=28
M296 1734 170 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.46824e-13 pd=8e-07 ps=1.22353e-06 nrd=0.166667 nrs=0.407843 sa=7.24e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=56340 $Y=32290 $D=28
M297 209 1733 1734 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=1.044e-06 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=56660 $Y=32290 $D=28
M298 1735 1733 209 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.524e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=57140 $Y=32290 $D=28
M299 VSS 170 1735 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=1.844e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=57460 $Y=32290 $D=28
M300 VSS 246 1736 VSS lpnfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02776e-13 as=1.344e-13 pd=8.56471e-07 ps=1.48e-06 nrd=0.582633 nrs=0.761905 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=65780 $Y=56090 $D=28
M301 1737 241 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.46824e-13 pd=8e-07 ps=1.22353e-06 nrd=0.166667 nrs=0.407843 sa=7.24e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=66340 $Y=55910 $D=28
M302 247 1736 1737 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=1.044e-06 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=66660 $Y=55910 $D=28
M303 1738 1736 247 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.524e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=67140 $Y=55910 $D=28
M304 VSS 241 1738 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=1.844e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=67460 $Y=55910 $D=28
M305 VSS 742 1739 VSS lpnfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02776e-13 as=1.344e-13 pd=8.56471e-07 ps=1.48e-06 nrd=0.582633 nrs=0.761905 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=186180 $Y=53890 $D=28
M306 1740 788 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.46824e-13 pd=8e-07 ps=1.22353e-06 nrd=0.166667 nrs=0.407843 sa=7.24e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=186740 $Y=53890 $D=28
M307 869 1739 1740 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=1.044e-06 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=187060 $Y=53890 $D=28
M308 1741 1739 869 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.524e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=187540 $Y=53890 $D=28
M309 VSS 788 1741 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=1.844e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=187860 $Y=53890 $D=28
M310 VSS 55 1742 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.17727e-13 as=1.408e-13 pd=8.74634e-07 ps=1.52e-06 nrd=0.608093 nrs=0.727273 sa=3.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=14880 $Y=70450 $D=28
M311 37 1742 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.46156e-13 pd=1.28e-06 ps=1.82878e-06 nrd=0.195652 nrs=0.290827 sa=6.05217e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=15440 $Y=69990 $D=28
M312 VSS 23 37 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.08522e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=15920 $Y=69990 $D=28
M313 VSS 101 1745 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.17727e-13 as=1.408e-13 pd=8.74634e-07 ps=1.52e-06 nrd=0.608093 nrs=0.727273 sa=3.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=27280 $Y=32310 $D=28
M314 52 1745 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.46156e-13 pd=1.28e-06 ps=1.82878e-06 nrd=0.195652 nrs=0.290827 sa=6.05217e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=27840 $Y=32290 $D=28
M315 VSS 199 52 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.08522e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=28320 $Y=32290 $D=28
M316 VSS 129 1748 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.17727e-13 as=1.408e-13 pd=8.74634e-07 ps=1.52e-06 nrd=0.608093 nrs=0.727273 sa=3.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=37680 $Y=41650 $D=28
M317 140 1748 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.46156e-13 pd=1.28e-06 ps=1.82878e-06 nrd=0.195652 nrs=0.290827 sa=6.05217e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=38240 $Y=41190 $D=28
M318 VSS 82 140 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.08522e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=38720 $Y=41190 $D=28
M319 VSS 394 1751 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.17727e-13 as=1.408e-13 pd=8.74634e-07 ps=1.52e-06 nrd=0.608093 nrs=0.727273 sa=3.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=100880 $Y=56050 $D=28
M320 369 1751 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.46156e-13 pd=1.28e-06 ps=1.82878e-06 nrd=0.195652 nrs=0.290827 sa=6.05217e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=101440 $Y=55590 $D=28
M321 VSS 437 369 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.08522e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=101920 $Y=55590 $D=28
M322 VSS 913 1754 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.17727e-13 as=1.408e-13 pd=8.74634e-07 ps=1.52e-06 nrd=0.608093 nrs=0.727273 sa=3.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=141280 $Y=68310 $D=28
M323 552 1754 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.46156e-13 pd=1.28e-06 ps=1.82878e-06 nrd=0.195652 nrs=0.290827 sa=6.05217e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=141840 $Y=68290 $D=28
M324 VSS 561 552 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.08522e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=142320 $Y=68290 $D=28
M325 VSS 868 1757 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.17727e-13 as=1.408e-13 pd=8.74634e-07 ps=1.52e-06 nrd=0.608093 nrs=0.727273 sa=3.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=186480 $Y=34450 $D=28
M326 781 1757 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.46156e-13 pd=1.28e-06 ps=1.82878e-06 nrd=0.195652 nrs=0.290827 sa=6.05217e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=187040 $Y=33990 $D=28
M327 VSS 771 781 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.08522e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=187520 $Y=33990 $D=28
M328 VSS 869 1760 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.17727e-13 as=1.408e-13 pd=8.74634e-07 ps=1.52e-06 nrd=0.608093 nrs=0.727273 sa=3.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=186480 $Y=41650 $D=28
M329 782 1760 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.46156e-13 pd=1.28e-06 ps=1.82878e-06 nrd=0.195652 nrs=0.290827 sa=6.05217e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=187040 $Y=41190 $D=28
M330 VSS 779 782 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.08522e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=187520 $Y=41190 $D=28
M331 1764 21 1763 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.44e-14 pd=4e-07 ps=1.28e-06 nrd=0.5 nrs=2.36 sa=3.6e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=8960 $Y=34590 $D=28
M332 VSS 17 1764 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92708e-14 as=2e-14 pd=6.83333e-07 ps=4e-07 nrd=1.98177 nrs=0.5 sa=6.8e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=9280 $Y=34590 $D=28
M333 38 1763 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.9025e-13 pd=1.6e-06 ps=1.64e-06 nrd=0.666667 nrs=0.825738 sa=7.20833e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=9840 $Y=34430 $D=28
M334 1766 825 1765 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.44e-14 pd=4e-07 ps=1.28e-06 nrd=0.5 nrs=2.36 sa=3.6e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=75360 $Y=25210 $D=28
M335 VSS 281 1766 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92708e-14 as=2e-14 pd=6.83333e-07 ps=4e-07 nrd=1.98177 nrs=0.5 sa=6.8e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=75680 $Y=25210 $D=28
M336 826 1765 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.9025e-13 pd=1.6e-06 ps=1.64e-06 nrd=0.666667 nrs=0.825738 sa=7.20833e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=76240 $Y=25090 $D=28
M337 1768 525 1767 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.44e-14 pd=4e-07 ps=1.28e-06 nrd=0.5 nrs=2.36 sa=3.6e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=129360 $Y=46810 $D=28
M338 VSS 517 1768 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92708e-14 as=2e-14 pd=6.83333e-07 ps=4e-07 nrd=1.98177 nrs=0.5 sa=6.8e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=129680 $Y=46810 $D=28
M339 498 1767 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.9025e-13 pd=1.6e-06 ps=1.64e-06 nrd=0.666667 nrs=0.825738 sa=7.20833e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=130240 $Y=46690 $D=28
M340 1770 501 1769 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.44e-14 pd=4e-07 ps=1.28e-06 nrd=0.5 nrs=2.36 sa=3.6e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=130960 $Y=27390 $D=28
M341 VSS 504 1770 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92708e-14 as=2e-14 pd=6.83333e-07 ps=4e-07 nrd=1.98177 nrs=0.5 sa=6.8e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=131280 $Y=27390 $D=28
M342 507 1769 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.9025e-13 pd=1.6e-06 ps=1.64e-06 nrd=0.666667 nrs=0.825738 sa=7.20833e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=131840 $Y=27230 $D=28
M343 1772 558 1771 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.44e-14 pd=4e-07 ps=1.28e-06 nrd=0.5 nrs=2.36 sa=3.6e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=143760 $Y=32410 $D=28
M344 VSS 554 1772 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92708e-14 as=2e-14 pd=6.83333e-07 ps=4e-07 nrd=1.98177 nrs=0.5 sa=6.8e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=144080 $Y=32410 $D=28
M345 573 1771 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.9025e-13 pd=1.6e-06 ps=1.64e-06 nrd=0.666667 nrs=0.825738 sa=7.20833e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=144640 $Y=32290 $D=28
M346 1774 642 1773 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.44e-14 pd=4e-07 ps=1.28e-06 nrd=0.5 nrs=2.36 sa=3.6e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=159360 $Y=48990 $D=28
M347 VSS 633 1774 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92708e-14 as=2e-14 pd=6.83333e-07 ps=4e-07 nrd=1.98177 nrs=0.5 sa=6.8e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=159680 $Y=48990 $D=28
M348 634 1773 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.9025e-13 pd=1.6e-06 ps=1.64e-06 nrd=0.666667 nrs=0.825738 sa=7.20833e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=160240 $Y=48830 $D=28
M349 1776 625 1775 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.44e-14 pd=4e-07 ps=1.28e-06 nrd=0.5 nrs=2.36 sa=3.6e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=164560 $Y=46810 $D=28
M350 VSS 660 1776 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92708e-14 as=2e-14 pd=6.83333e-07 ps=4e-07 nrd=1.98177 nrs=0.5 sa=6.8e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=164880 $Y=46810 $D=28
M351 663 1775 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.9025e-13 pd=1.6e-06 ps=1.64e-06 nrd=0.666667 nrs=0.825738 sa=7.20833e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=165440 $Y=46690 $D=28
M352 1778 677 1777 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.44e-14 pd=4e-07 ps=1.28e-06 nrd=0.5 nrs=2.36 sa=3.6e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=166160 $Y=68410 $D=28
M353 VSS 692 1778 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92708e-14 as=2e-14 pd=6.83333e-07 ps=4e-07 nrd=1.98177 nrs=0.5 sa=6.8e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=166480 $Y=68410 $D=28
M354 672 1777 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.9025e-13 pd=1.6e-06 ps=1.64e-06 nrd=0.666667 nrs=0.825738 sa=7.20833e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=167040 $Y=68290 $D=28
M355 1780 684 1779 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.44e-14 pd=4e-07 ps=1.28e-06 nrd=0.5 nrs=2.36 sa=3.6e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=168160 $Y=63390 $D=28
M356 VSS 679 1780 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92708e-14 as=2e-14 pd=6.83333e-07 ps=4e-07 nrd=1.98177 nrs=0.5 sa=6.8e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=168480 $Y=63390 $D=28
M357 861 1779 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.9025e-13 pd=1.6e-06 ps=1.64e-06 nrd=0.666667 nrs=0.825738 sa=7.20833e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=169040 $Y=63230 $D=28
M358 1782 707 1781 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.44e-14 pd=4e-07 ps=1.28e-06 nrd=0.5 nrs=2.36 sa=3.6e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=177360 $Y=63390 $D=28
M359 VSS 736 1782 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92708e-14 as=2e-14 pd=6.83333e-07 ps=4e-07 nrd=1.98177 nrs=0.5 sa=6.8e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=177680 $Y=63390 $D=28
M360 738 1781 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.9025e-13 pd=1.6e-06 ps=1.64e-06 nrd=0.666667 nrs=0.825738 sa=7.20833e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=178240 $Y=63230 $D=28
M361 1784 778 1783 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.44e-14 pd=4e-07 ps=1.28e-06 nrd=0.5 nrs=2.36 sa=3.6e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=179360 $Y=41790 $D=28
M362 VSS 757 1784 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92708e-14 as=2e-14 pd=6.83333e-07 ps=4e-07 nrd=1.98177 nrs=0.5 sa=6.8e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=179680 $Y=41790 $D=28
M363 749 1783 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.9025e-13 pd=1.6e-06 ps=1.64e-06 nrd=0.666667 nrs=0.825738 sa=7.20833e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=180240 $Y=41630 $D=28
M364 1786 770 1785 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.44e-14 pd=4e-07 ps=1.28e-06 nrd=0.5 nrs=2.36 sa=3.6e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=184960 $Y=18010 $D=28
M365 VSS 772 1786 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92708e-14 as=2e-14 pd=6.83333e-07 ps=4e-07 nrd=1.98177 nrs=0.5 sa=6.8e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=185280 $Y=18010 $D=28
M366 774 1785 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.9025e-13 pd=1.6e-06 ps=1.64e-06 nrd=0.666667 nrs=0.825738 sa=7.20833e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=185840 $Y=17890 $D=28
M367 43 124 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=18860 $Y=53890 $D=28
M368 VSS 44 43 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=19340 $Y=53890 $D=28
M369 65 81 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=21660 $Y=68290 $D=28
M370 VSS 80 65 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=22140 $Y=68290 $D=28
M371 146 107 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=42860 $Y=48390 $D=28
M372 VSS 98 146 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=43340 $Y=48390 $D=28
M373 156 131 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=44860 $Y=48390 $D=28
M374 VSS 82 156 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=45340 $Y=48390 $D=28
M375 249 244 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=67260 $Y=25090 $D=28
M376 VSS 243 249 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=67740 $Y=25090 $D=28
M377 357 378 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=106060 $Y=41190 $D=28
M378 VSS 409 357 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=106540 $Y=41190 $D=28
M379 442 431 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=116060 $Y=75490 $D=28
M380 VSS 439 442 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=116540 $Y=75490 $D=28
M381 497 480 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=126860 $Y=39490 $D=28
M382 VSS 845 497 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=127340 $Y=39490 $D=28
M383 494 487 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=128460 $Y=55590 $D=28
M384 VSS 485 494 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=128940 $Y=55590 $D=28
M385 492 470 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=132860 $Y=41190 $D=28
M386 VSS 493 492 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=133340 $Y=41190 $D=28
M387 852 514 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=133660 $Y=19590 $D=28
M388 VSS 491 852 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=134140 $Y=19590 $D=28
M389 540 535 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=137660 $Y=39490 $D=28
M390 VSS 500 540 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=138140 $Y=39490 $D=28
M391 669 497 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=139660 $Y=46690 $D=28
M392 VSS 512 669 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=140140 $Y=46690 $D=28
M393 856 590 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=145660 $Y=68290 $D=28
M394 VSS 575 856 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=146140 $Y=68290 $D=28
M395 858 705 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=156860 $Y=68290 $D=28
M396 VSS 575 858 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=157340 $Y=68290 $D=28
M397 636 667 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=162460 $Y=55590 $D=28
M398 VSS 648 636 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=162940 $Y=55590 $D=28
M399 859 644 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=166060 $Y=75490 $D=28
M400 VSS 575 859 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=166540 $Y=75490 $D=28
M401 754 767 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=180460 $Y=17890 $D=28
M402 VSS 693 754 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=180940 $Y=17890 $D=28
M403 762 777 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=182060 $Y=61090 $D=28
M404 VSS 681 762 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=182540 $Y=61090 $D=28
M405 864 768 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.916e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.344518 sa=3.16957e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=184460 $Y=41190 $D=28
M406 VSS 681 864 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=7.96957e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=184940 $Y=41190 $D=28
M407 1828 15 63 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=9360 $Y=19590 $D=28
M408 VSS 29 1828 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=9680 $Y=19590 $D=28
M409 1829 29 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=10280 $Y=19590 $D=28
M410 63 15 1829 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=10600 $Y=19590 $D=28
M411 1830 15 63 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=11080 $Y=19590 $D=28
M412 VSS 29 1830 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=11400 $Y=19590 $D=28
M413 63 799 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=12020 $Y=19590 $D=28
M414 VSS 799 63 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=12500 $Y=19900 $D=28
M415 63 799 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=12980 $Y=19900 $D=28
M416 1832 207 118 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=52160 $Y=17990 $D=28
M417 VSS 235 1832 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=52480 $Y=17990 $D=28
M418 1833 235 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=53080 $Y=17990 $D=28
M419 118 207 1833 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=53400 $Y=17990 $D=28
M420 1834 207 118 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=53880 $Y=17990 $D=28
M421 VSS 235 1834 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=54200 $Y=17990 $D=28
M422 118 208 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=54820 $Y=17990 $D=28
M423 VSS 208 118 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=55300 $Y=17990 $D=28
M424 118 208 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=55780 $Y=17990 $D=28
M425 1836 405 834 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=108160 $Y=32390 $D=28
M426 VSS 445 1836 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=108480 $Y=32390 $D=28
M427 1837 445 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=109080 $Y=32390 $D=28
M428 834 405 1837 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=109400 $Y=32390 $D=28
M429 1838 405 834 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=109880 $Y=32390 $D=28
M430 VSS 445 1838 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=110200 $Y=32390 $D=28
M431 834 409 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=110820 $Y=32390 $D=28
M432 VSS 409 834 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=111300 $Y=32390 $D=28
M433 834 409 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=111780 $Y=32390 $D=28
M434 1840 467 495 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=120560 $Y=62790 $D=28
M435 VSS 460 1840 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=120880 $Y=62790 $D=28
M436 1841 460 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=121480 $Y=62790 $D=28
M437 495 467 1841 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=121800 $Y=62790 $D=28
M438 1842 467 495 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=122280 $Y=62790 $D=28
M439 VSS 460 1842 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=122600 $Y=62790 $D=28
M440 495 462 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=123220 $Y=62790 $D=28
M441 VSS 462 495 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=123700 $Y=63100 $D=28
M442 495 462 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=124180 $Y=63100 $D=28
M443 1844 545 441 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=121760 $Y=39590 $D=28
M444 VSS 488 1844 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=122080 $Y=39590 $D=28
M445 1845 488 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=122680 $Y=39590 $D=28
M446 441 545 1845 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=123000 $Y=39590 $D=28
M447 1846 545 441 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=123480 $Y=39590 $D=28
M448 VSS 488 1846 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=123800 $Y=39590 $D=28
M449 441 506 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=124420 $Y=39590 $D=28
M450 VSS 506 441 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=124900 $Y=39590 $D=28
M451 441 506 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=125380 $Y=39590 $D=28
M452 1848 404 842 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=121760 $Y=75590 $D=28
M453 VSS 490 1848 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=122080 $Y=75590 $D=28
M454 1849 490 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=122680 $Y=75590 $D=28
M455 842 404 1849 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=123000 $Y=75590 $D=28
M456 1850 404 842 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=123480 $Y=75590 $D=28
M457 VSS 490 1850 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=123800 $Y=75590 $D=28
M458 842 482 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=124420 $Y=75590 $D=28
M459 VSS 482 842 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=124900 $Y=75590 $D=28
M460 842 482 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=125380 $Y=75590 $D=28
M461 1852 499 483 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=124160 $Y=32390 $D=28
M462 VSS 472 1852 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=124480 $Y=32390 $D=28
M463 1853 472 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=125080 $Y=32390 $D=28
M464 483 499 1853 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=125400 $Y=32390 $D=28
M465 1854 499 483 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=125880 $Y=32390 $D=28
M466 VSS 472 1854 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=126200 $Y=32390 $D=28
M467 483 459 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=126820 $Y=32390 $D=28
M468 VSS 459 483 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=127300 $Y=32390 $D=28
M469 483 459 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=127780 $Y=32390 $D=28
M470 1856 499 571 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=132560 $Y=33990 $D=28
M471 VSS 516 1856 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=132880 $Y=33990 $D=28
M472 1857 516 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=133480 $Y=33990 $D=28
M473 571 499 1857 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=133800 $Y=33990 $D=28
M474 1858 499 571 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=134280 $Y=33990 $D=28
M475 VSS 516 1858 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=134600 $Y=33990 $D=28
M476 571 537 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=135220 $Y=33990 $D=28
M477 VSS 537 571 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=135700 $Y=34300 $D=28
M478 571 537 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=136180 $Y=34300 $D=28
M479 1860 545 542 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=139360 $Y=39590 $D=28
M480 VSS 547 1860 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=139680 $Y=39590 $D=28
M481 1861 547 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=140280 $Y=39590 $D=28
M482 542 545 1861 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=140600 $Y=39590 $D=28
M483 1862 545 542 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=141080 $Y=39590 $D=28
M484 VSS 547 1862 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=141400 $Y=39590 $D=28
M485 542 531 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=142020 $Y=39590 $D=28
M486 VSS 531 542 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=142500 $Y=39590 $D=28
M487 542 531 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=142980 $Y=39590 $D=28
M488 1864 545 583 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=139360 $Y=55590 $D=28
M489 VSS 565 1864 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=139680 $Y=55590 $D=28
M490 1865 565 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=140280 $Y=55590 $D=28
M491 583 545 1865 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=140600 $Y=55590 $D=28
M492 1866 545 583 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=141080 $Y=55590 $D=28
M493 VSS 565 1866 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=141400 $Y=55590 $D=28
M494 583 572 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=142020 $Y=55590 $D=28
M495 VSS 572 583 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=142500 $Y=55900 $D=28
M496 583 572 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=142980 $Y=55900 $D=28
M497 1868 562 702 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=169360 $Y=48390 $D=28
M498 VSS 691 1868 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=169680 $Y=48390 $D=28
M499 1869 691 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=170280 $Y=48390 $D=28
M500 702 562 1869 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=170600 $Y=48390 $D=28
M501 1870 562 702 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=171080 $Y=48390 $D=28
M502 VSS 691 1870 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=171400 $Y=48390 $D=28
M503 702 739 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=172020 $Y=48390 $D=28
M504 VSS 739 702 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=172500 $Y=48700 $D=28
M505 702 739 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=172980 $Y=48700 $D=28
M506 1872 742 764 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=176560 $Y=32390 $D=28
M507 VSS 737 1872 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=176880 $Y=32390 $D=28
M508 1873 737 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=177480 $Y=32390 $D=28
M509 764 742 1873 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=177800 $Y=32390 $D=28
M510 1874 742 764 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=178280 $Y=32390 $D=28
M511 VSS 737 1874 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=178600 $Y=32390 $D=28
M512 764 741 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=179220 $Y=32390 $D=28
M513 VSS 741 764 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=179700 $Y=32390 $D=28
M514 764 741 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=180180 $Y=32390 $D=28
M515 1876 729 751 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=176960 $Y=61190 $D=28
M516 VSS 776 1876 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=177280 $Y=61190 $D=28
M517 1877 776 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=177880 $Y=61190 $D=28
M518 751 729 1877 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=178200 $Y=61190 $D=28
M519 1878 729 751 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=178680 $Y=61190 $D=28
M520 VSS 776 1878 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=179000 $Y=61190 $D=28
M521 751 786 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=179620 $Y=61190 $D=28
M522 VSS 786 751 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=180100 $Y=61190 $D=28
M523 751 786 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=180580 $Y=61190 $D=28
M524 1880 729 763 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=179360 $Y=69990 $D=28
M525 VSS 745 1880 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=179680 $Y=69990 $D=28
M526 1881 745 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=180280 $Y=69990 $D=28
M527 763 729 1881 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=180600 $Y=69990 $D=28
M528 1882 729 763 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=181080 $Y=69990 $D=28
M529 VSS 745 1882 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=181400 $Y=69990 $D=28
M530 763 758 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=182020 $Y=69990 $D=28
M531 VSS 758 763 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=182500 $Y=70300 $D=28
M532 763 758 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=182980 $Y=70300 $D=28
M533 1884 755 787 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=2.624e-13 pd=1.02e-06 ps=2.28e-06 nrd=0.121951 nrs=0.390244 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=184160 $Y=25190 $D=28
M534 VSS 742 1884 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.968e-13 as=8.2e-14 pd=1.3e-06 ps=1.02e-06 nrd=0.292683 nrs=0.121951 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=184480 $Y=25190 $D=28
M535 1885 742 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.968e-13 pd=1.02e-06 ps=1.3e-06 nrd=0.121951 nrs=0.292683 sa=1.24e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=185080 $Y=25190 $D=28
M536 787 755 1885 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.56e-06 sb=1.88659e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=185400 $Y=25190 $D=28
M537 1886 755 787 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=1.70512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=185880 $Y=25190 $D=28
M538 VSS 742 1886 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.05e-13 as=8.2e-14 pd=1.32e-06 ps=1.02e-06 nrd=0.304878 nrs=0.121951 sa=2e-06 sb=1.52195e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=186200 $Y=25190 $D=28
M539 787 780 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66713e-13 as=2.05e-13 pd=1.45504e-06 ps=1.32e-06 nrd=0.247937 nrs=0.304878 sa=2e-06 sb=9.01951e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=186820 $Y=25190 $D=28
M540 VSS 780 787 VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.18e-14 as=1.03687e-13 pd=8.7e-07 ps=9.04962e-07 nrd=0.352941 nrs=0.398644 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=187300 $Y=25190 $D=28
M541 787 780 VSS VSS lpnfet w=5.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.632e-13 as=9.18e-14 pd=1.66e-06 ps=8.7e-07 nrd=0.627451 nrs=0.352941 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=187780 $Y=25190 $D=28
M542 1888 411 383 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.92e-13 pd=8e-07 ps=1.84e-06 nrd=0.166667 nrs=0.533333 sa=3.2e-07 sb=1.872e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=104800 $Y=75490 $D=28
M543 VSS 387 1888 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.74e-13 as=6e-14 pd=1.32162e-06 ps=8e-07 nrd=0.483333 nrs=0.166667 sa=6.4e-07 sb=1.79733e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=105120 $Y=75490 $D=28
M544 1889 387 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.74e-13 pd=8e-07 ps=1.32162e-06 nrd=0.166667 nrs=0.483333 sa=1.2e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=105680 $Y=75490 $D=28
M545 383 411 1889 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.1366e-13 as=6e-14 pd=1.08679e-06 ps=8e-07 nrd=0.315723 nrs=0.166667 sa=1.52e-06 sb=1.04e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=106000 $Y=75490 $D=28
M546 VSS 393 383 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=8.71396e-14 pd=8.2e-07 ps=8.33208e-07 nrd=0.391304 nrs=0.411813 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=106480 $Y=75540 $D=28
M547 383 393 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=8.28e-14 pd=1.56e-06 ps=8.2e-07 nrd=0.695652 nrs=0.391304 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=106960 $Y=75540 $D=28
M548 1891 422 833 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.92e-13 pd=8e-07 ps=1.84e-06 nrd=0.166667 nrs=0.533333 sa=3.2e-07 sb=1.872e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=108800 $Y=63110 $D=28
M549 VSS 411 1891 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.74e-13 as=6e-14 pd=1.32162e-06 ps=8e-07 nrd=0.483333 nrs=0.166667 sa=6.4e-07 sb=1.79733e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=109120 $Y=63110 $D=28
M550 1892 411 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.74e-13 pd=8e-07 ps=1.32162e-06 nrd=0.166667 nrs=0.483333 sa=1.2e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=109680 $Y=63110 $D=28
M551 833 422 1892 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.1366e-13 as=6e-14 pd=1.08679e-06 ps=8e-07 nrd=0.315723 nrs=0.166667 sa=1.52e-06 sb=1.04e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=110000 $Y=63110 $D=28
M552 VSS 420 833 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=8.71396e-14 pd=8.2e-07 ps=8.33208e-07 nrd=0.391304 nrs=0.411813 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=110480 $Y=63200 $D=28
M553 833 420 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=8.28e-14 pd=1.56e-06 ps=8.2e-07 nrd=0.695652 nrs=0.391304 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=110960 $Y=63200 $D=28
M554 1894 411 464 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.92e-13 pd=8e-07 ps=1.84e-06 nrd=0.166667 nrs=0.533333 sa=3.2e-07 sb=1.872e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=118000 $Y=75490 $D=28
M555 VSS 442 1894 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.74e-13 as=6e-14 pd=1.32162e-06 ps=8e-07 nrd=0.483333 nrs=0.166667 sa=6.4e-07 sb=1.79733e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=118320 $Y=75490 $D=28
M556 1895 442 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.74e-13 pd=8e-07 ps=1.32162e-06 nrd=0.166667 nrs=0.483333 sa=1.2e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=118880 $Y=75490 $D=28
M557 464 411 1895 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.1366e-13 as=6e-14 pd=1.08679e-06 ps=8e-07 nrd=0.315723 nrs=0.166667 sa=1.52e-06 sb=1.04e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=119200 $Y=75490 $D=28
M558 VSS 840 464 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=8.71396e-14 pd=8.2e-07 ps=8.33208e-07 nrd=0.391304 nrs=0.411813 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=119680 $Y=75540 $D=28
M559 464 840 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=8.28e-14 pd=1.56e-06 ps=8.2e-07 nrd=0.695652 nrs=0.391304 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=120160 $Y=75540 $D=28
M560 1897 518 511 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.92e-13 pd=8e-07 ps=1.84e-06 nrd=0.166667 nrs=0.533333 sa=3.2e-07 sb=1.872e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=133600 $Y=55910 $D=28
M561 VSS 524 1897 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.74e-13 as=6e-14 pd=1.32162e-06 ps=8e-07 nrd=0.483333 nrs=0.166667 sa=6.4e-07 sb=1.79733e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=133920 $Y=55910 $D=28
M562 1898 524 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.74e-13 pd=8e-07 ps=1.32162e-06 nrd=0.166667 nrs=0.483333 sa=1.2e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=134480 $Y=55910 $D=28
M563 511 518 1898 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.1366e-13 as=6e-14 pd=1.08679e-06 ps=8e-07 nrd=0.315723 nrs=0.166667 sa=1.52e-06 sb=1.04e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=134800 $Y=55910 $D=28
M564 VSS 534 511 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=8.71396e-14 pd=8.2e-07 ps=8.33208e-07 nrd=0.391304 nrs=0.411813 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=135280 $Y=56000 $D=28
M565 511 534 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=8.28e-14 pd=1.56e-06 ps=8.2e-07 nrd=0.695652 nrs=0.391304 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=135760 $Y=56000 $D=28
M566 1900 912 532 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.92e-13 pd=8e-07 ps=1.84e-06 nrd=0.166667 nrs=0.533333 sa=3.2e-07 sb=1.872e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=137200 $Y=41510 $D=28
M567 VSS 510 1900 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.74e-13 as=6e-14 pd=1.32162e-06 ps=8e-07 nrd=0.483333 nrs=0.166667 sa=6.4e-07 sb=1.79733e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=137520 $Y=41510 $D=28
M568 1901 510 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.74e-13 pd=8e-07 ps=1.32162e-06 nrd=0.166667 nrs=0.483333 sa=1.2e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=138080 $Y=41510 $D=28
M569 532 912 1901 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.1366e-13 as=6e-14 pd=1.08679e-06 ps=8e-07 nrd=0.315723 nrs=0.166667 sa=1.52e-06 sb=1.04e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=138400 $Y=41510 $D=28
M570 VSS 546 532 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=8.71396e-14 pd=8.2e-07 ps=8.33208e-07 nrd=0.391304 nrs=0.411813 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=138880 $Y=41600 $D=28
M571 532 546 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=8.28e-14 pd=1.56e-06 ps=8.2e-07 nrd=0.695652 nrs=0.391304 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=139360 $Y=41600 $D=28
M572 1903 594 587 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.92e-13 pd=8e-07 ps=1.84e-06 nrd=0.166667 nrs=0.533333 sa=3.2e-07 sb=1.872e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=150400 $Y=48710 $D=28
M573 VSS 669 1903 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.74e-13 as=6e-14 pd=1.32162e-06 ps=8e-07 nrd=0.483333 nrs=0.166667 sa=6.4e-07 sb=1.79733e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=150720 $Y=48710 $D=28
M574 1904 669 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.74e-13 pd=8e-07 ps=1.32162e-06 nrd=0.166667 nrs=0.483333 sa=1.2e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=151280 $Y=48710 $D=28
M575 587 594 1904 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.1366e-13 as=6e-14 pd=1.08679e-06 ps=8e-07 nrd=0.315723 nrs=0.166667 sa=1.52e-06 sb=1.04e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=151600 $Y=48710 $D=28
M576 VSS 598 587 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=8.71396e-14 pd=8.2e-07 ps=8.33208e-07 nrd=0.391304 nrs=0.411813 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=152080 $Y=48800 $D=28
M577 587 598 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=8.28e-14 pd=1.56e-06 ps=8.2e-07 nrd=0.695652 nrs=0.391304 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=152560 $Y=48800 $D=28
M578 1906 562 857 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.92e-13 pd=8e-07 ps=1.84e-06 nrd=0.166667 nrs=0.533333 sa=3.2e-07 sb=1.872e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=158800 $Y=68290 $D=28
M579 VSS 636 1906 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.74e-13 as=6e-14 pd=1.32162e-06 ps=8e-07 nrd=0.483333 nrs=0.166667 sa=6.4e-07 sb=1.79733e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=159120 $Y=68290 $D=28
M580 1907 636 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.74e-13 pd=8e-07 ps=1.32162e-06 nrd=0.166667 nrs=0.483333 sa=1.2e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=159680 $Y=68290 $D=28
M581 857 562 1907 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.1366e-13 as=6e-14 pd=1.08679e-06 ps=8e-07 nrd=0.315723 nrs=0.166667 sa=1.52e-06 sb=1.04e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=160000 $Y=68290 $D=28
M582 VSS 674 857 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=8.71396e-14 pd=8.2e-07 ps=8.33208e-07 nrd=0.391304 nrs=0.411813 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=160480 $Y=68340 $D=28
M583 857 674 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=8.28e-14 pd=1.56e-06 ps=8.2e-07 nrd=0.695652 nrs=0.391304 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=160960 $Y=68340 $D=28
M584 1909 518 637 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.92e-13 pd=8e-07 ps=1.84e-06 nrd=0.166667 nrs=0.533333 sa=3.2e-07 sb=1.872e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=159600 $Y=53890 $D=28
M585 VSS 653 1909 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.74e-13 as=6e-14 pd=1.32162e-06 ps=8e-07 nrd=0.483333 nrs=0.166667 sa=6.4e-07 sb=1.79733e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=159920 $Y=53890 $D=28
M586 1910 653 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.74e-13 pd=8e-07 ps=1.32162e-06 nrd=0.166667 nrs=0.483333 sa=1.2e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=160480 $Y=53890 $D=28
M587 637 518 1910 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.1366e-13 as=6e-14 pd=1.08679e-06 ps=8e-07 nrd=0.315723 nrs=0.166667 sa=1.52e-06 sb=1.04e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=160800 $Y=53890 $D=28
M588 VSS 650 637 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=8.71396e-14 pd=8.2e-07 ps=8.33208e-07 nrd=0.391304 nrs=0.411813 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=161280 $Y=53940 $D=28
M589 637 650 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=8.28e-14 pd=1.56e-06 ps=8.2e-07 nrd=0.695652 nrs=0.391304 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=161760 $Y=53940 $D=28
M590 1912 598 690 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.92e-13 pd=8e-07 ps=1.84e-06 nrd=0.166667 nrs=0.533333 sa=3.2e-07 sb=1.872e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=166000 $Y=48710 $D=28
M591 VSS 710 1912 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.74e-13 as=6e-14 pd=1.32162e-06 ps=8e-07 nrd=0.483333 nrs=0.166667 sa=6.4e-07 sb=1.79733e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=166320 $Y=48710 $D=28
M592 1913 710 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.74e-13 pd=8e-07 ps=1.32162e-06 nrd=0.166667 nrs=0.483333 sa=1.2e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=166880 $Y=48710 $D=28
M593 690 598 1913 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.1366e-13 as=6e-14 pd=1.08679e-06 ps=8e-07 nrd=0.315723 nrs=0.166667 sa=1.52e-06 sb=1.04e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=167200 $Y=48710 $D=28
M594 VSS 727 690 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=8.71396e-14 pd=8.2e-07 ps=8.33208e-07 nrd=0.391304 nrs=0.411813 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=167680 $Y=48800 $D=28
M595 690 727 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=8.28e-14 pd=1.56e-06 ps=8.2e-07 nrd=0.695652 nrs=0.391304 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=168160 $Y=48800 $D=28
M596 1915 674 784 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.92e-13 pd=8e-07 ps=1.84e-06 nrd=0.166667 nrs=0.533333 sa=3.2e-07 sb=1.872e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=168000 $Y=61090 $D=28
M597 VSS 696 1915 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.74e-13 as=6e-14 pd=1.32162e-06 ps=8e-07 nrd=0.483333 nrs=0.166667 sa=6.4e-07 sb=1.79733e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=168320 $Y=61090 $D=28
M598 1916 696 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.74e-13 pd=8e-07 ps=1.32162e-06 nrd=0.166667 nrs=0.483333 sa=1.2e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=168880 $Y=61090 $D=28
M599 784 674 1916 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.1366e-13 as=6e-14 pd=1.08679e-06 ps=8e-07 nrd=0.315723 nrs=0.166667 sa=1.52e-06 sb=1.04e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=169200 $Y=61090 $D=28
M600 VSS 728 784 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=8.71396e-14 pd=8.2e-07 ps=8.33208e-07 nrd=0.391304 nrs=0.411813 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=169680 $Y=61140 $D=28
M601 784 728 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=8.28e-14 pd=1.56e-06 ps=8.2e-07 nrd=0.695652 nrs=0.391304 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=170160 $Y=61140 $D=28
M602 1918 518 866 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.92e-13 pd=8e-07 ps=1.84e-06 nrd=0.166667 nrs=0.533333 sa=3.2e-07 sb=1.872e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=184000 $Y=61090 $D=28
M603 VSS 769 1918 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.74e-13 as=6e-14 pd=1.32162e-06 ps=8e-07 nrd=0.483333 nrs=0.166667 sa=6.4e-07 sb=1.79733e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=184320 $Y=61090 $D=28
M604 1919 769 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.74e-13 pd=8e-07 ps=1.32162e-06 nrd=0.166667 nrs=0.483333 sa=1.2e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=184880 $Y=61090 $D=28
M605 866 518 1919 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.1366e-13 as=6e-14 pd=1.08679e-06 ps=8e-07 nrd=0.315723 nrs=0.166667 sa=1.52e-06 sb=1.04e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=185200 $Y=61090 $D=28
M606 VSS 775 866 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=8.71396e-14 pd=8.2e-07 ps=8.33208e-07 nrd=0.391304 nrs=0.411813 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=185680 $Y=61140 $D=28
M607 866 775 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=8.28e-14 pd=1.56e-06 ps=8.2e-07 nrd=0.695652 nrs=0.391304 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=186160 $Y=61140 $D=28
M608 1920 173 VSS VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92e-14 as=1.152e-13 pd=8e-07 ps=1.36e-06 nrd=0.611111 nrs=0.888889 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=47210 $Y=25250 $D=28
M609 VSS 140 1920 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.32846e-14 as=7.92e-14 pd=7.52308e-07 ps=8e-07 nrd=0.642628 nrs=0.611111 sa=8.8e-07 sb=7.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=47770 $Y=25250 $D=28
M610 147 1920 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.12838e-13 pd=2.48e-06 ps=1.92256e-06 nrd=0.347826 nrs=0.251463 sa=7.01413e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=48240 $Y=25090 $D=28
M611 1922 486 VSS VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92e-14 as=1.152e-13 pd=8e-07 ps=1.36e-06 nrd=0.611111 nrs=0.888889 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=123210 $Y=25250 $D=28
M612 VSS 474 1922 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.32846e-14 as=7.92e-14 pd=7.52308e-07 ps=8e-07 nrd=0.642628 nrs=0.611111 sa=8.8e-07 sb=7.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=123770 $Y=25250 $D=28
M613 501 1922 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.12838e-13 pd=2.48e-06 ps=1.92256e-06 nrd=0.347826 nrs=0.251463 sa=7.01413e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=124240 $Y=25090 $D=28
M614 1924 582 VSS VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92e-14 as=1.152e-13 pd=8e-07 ps=1.36e-06 nrd=0.611111 nrs=0.888889 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=147610 $Y=32450 $D=28
M615 VSS 573 1924 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.32846e-14 as=7.92e-14 pd=7.52308e-07 ps=8e-07 nrd=0.642628 nrs=0.611111 sa=8.8e-07 sb=7.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=148170 $Y=32450 $D=28
M616 591 1924 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.12838e-13 pd=2.48e-06 ps=1.92256e-06 nrd=0.347826 nrs=0.251463 sa=7.01413e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=148640 $Y=32290 $D=28
M617 1926 622 VSS VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92e-14 as=1.152e-13 pd=8e-07 ps=1.36e-06 nrd=0.611111 nrs=0.888889 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=154410 $Y=63190 $D=28
M618 VSS 609 1926 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.32846e-14 as=7.92e-14 pd=7.52308e-07 ps=8e-07 nrd=0.642628 nrs=0.611111 sa=8.8e-07 sb=7.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=154970 $Y=63190 $D=28
M619 602 1926 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.12838e-13 pd=2.48e-06 ps=1.92256e-06 nrd=0.347826 nrs=0.251463 sa=7.01413e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=155440 $Y=62790 $D=28
M620 1928 592 VSS VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92e-14 as=1.152e-13 pd=8e-07 ps=1.36e-06 nrd=0.611111 nrs=0.888889 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=155610 $Y=48790 $D=28
M621 VSS 634 1928 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.32846e-14 as=7.92e-14 pd=7.52308e-07 ps=8e-07 nrd=0.642628 nrs=0.611111 sa=8.8e-07 sb=7.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=156170 $Y=48790 $D=28
M622 600 1928 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.12838e-13 pd=2.48e-06 ps=1.92256e-06 nrd=0.347826 nrs=0.251463 sa=7.01413e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=156640 $Y=48390 $D=28
M623 1930 592 VSS VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92e-14 as=1.152e-13 pd=8e-07 ps=1.36e-06 nrd=0.611111 nrs=0.888889 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=157610 $Y=39650 $D=28
M624 VSS 663 1930 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.32846e-14 as=7.92e-14 pd=7.52308e-07 ps=8e-07 nrd=0.642628 nrs=0.611111 sa=8.8e-07 sb=7.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=158170 $Y=39650 $D=28
M625 574 1930 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.12838e-13 pd=2.48e-06 ps=1.92256e-06 nrd=0.347826 nrs=0.251463 sa=7.01413e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=158640 $Y=39490 $D=28
M626 1932 630 VSS VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92e-14 as=1.152e-13 pd=8e-07 ps=1.36e-06 nrd=0.611111 nrs=0.888889 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=158010 $Y=41590 $D=28
M627 VSS 646 1932 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.32846e-14 as=7.92e-14 pd=7.52308e-07 ps=8e-07 nrd=0.642628 nrs=0.611111 sa=8.8e-07 sb=7.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=158570 $Y=41590 $D=28
M628 625 1932 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.12838e-13 pd=2.48e-06 ps=1.92256e-06 nrd=0.347826 nrs=0.251463 sa=7.01413e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=159040 $Y=41190 $D=28
M629 1934 670 VSS VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92e-14 as=1.152e-13 pd=8e-07 ps=1.36e-06 nrd=0.611111 nrs=0.888889 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=164410 $Y=61250 $D=28
M630 VSS 576 1934 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.32846e-14 as=7.92e-14 pd=7.52308e-07 ps=8e-07 nrd=0.642628 nrs=0.611111 sa=8.8e-07 sb=7.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=164970 $Y=61250 $D=28
M631 684 1934 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.12838e-13 pd=2.48e-06 ps=1.92256e-06 nrd=0.347826 nrs=0.251463 sa=7.01413e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=165440 $Y=61090 $D=28
M632 1936 748 VSS VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92e-14 as=1.152e-13 pd=8e-07 ps=1.36e-06 nrd=0.611111 nrs=0.888889 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=182010 $Y=25250 $D=28
M633 VSS 717 1936 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.32846e-14 as=7.92e-14 pd=7.52308e-07 ps=8e-07 nrd=0.642628 nrs=0.611111 sa=8.8e-07 sb=7.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=182570 $Y=25250 $D=28
M634 761 1936 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.12838e-13 pd=2.48e-06 ps=1.92256e-06 nrd=0.347826 nrs=0.251463 sa=7.01413e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=183040 $Y=25090 $D=28
M635 1938 750 VSS VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.92e-14 as=1.152e-13 pd=8e-07 ps=1.36e-06 nrd=0.611111 nrs=0.888889 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=182810 $Y=54050 $D=28
M636 VSS 746 1938 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.32846e-14 as=7.92e-14 pd=7.52308e-07 ps=8e-07 nrd=0.642628 nrs=0.611111 sa=8.8e-07 sb=7.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=183370 $Y=54050 $D=28
M637 732 1938 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.12838e-13 pd=2.48e-06 ps=1.92256e-06 nrd=0.347826 nrs=0.251463 sa=7.01413e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=183840 $Y=53890 $D=28
M638 1940 52 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=12480 $Y=34310 $D=28
M639 34 70 1940 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=12800 $Y=34310 $D=28
M640 1941 40 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=14480 $Y=17890 $D=28
M641 19 29 1941 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=14800 $Y=17890 $D=28
M642 1942 30 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=15280 $Y=48710 $D=28
M643 35 14 1942 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=15600 $Y=48710 $D=28
M644 1943 36 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=16080 $Y=55910 $D=28
M645 31 48 1943 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=16400 $Y=55910 $D=28
M646 1944 44 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=17680 $Y=55910 $D=28
M647 36 124 1944 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=18000 $Y=55910 $D=28
M648 1945 44 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=20480 $Y=48710 $D=28
M649 61 124 1945 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=20800 $Y=48710 $D=28
M650 1946 91 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=20880 $Y=75490 $D=28
M651 64 67 1946 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=21200 $Y=75490 $D=28
M652 1947 132 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=37280 $Y=17890 $D=28
M653 116 137 1947 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=37600 $Y=17890 $D=28
M654 1948 140 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=45680 $Y=25090 $D=28
M655 154 173 1948 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=46000 $Y=25090 $D=28
M656 1949 198 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=54480 $Y=19910 $D=28
M657 243 814 1949 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=54800 $Y=19910 $D=28
M658 1950 815 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=58080 $Y=17890 $D=28
M659 816 207 1950 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=58400 $Y=17890 $D=28
M660 1951 243 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=65280 $Y=25090 $D=28
M661 258 244 1951 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=65600 $Y=25090 $D=28
M662 1952 258 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=70080 $Y=25090 $D=28
M663 259 262 1952 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=70400 $Y=25090 $D=28
M664 1953 904 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=70480 $Y=70310 $D=28
M665 277 289 1953 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=70800 $Y=70310 $D=28
M666 1954 274 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=73280 $Y=19910 $D=28
M667 281 298 1954 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=73600 $Y=19910 $D=28
M668 1955 297 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=76880 $Y=41510 $D=28
M669 292 286 1955 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=77200 $Y=41510 $D=28
M670 1956 361 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=96480 $Y=70310 $D=28
M671 909 830 1956 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=96800 $Y=70310 $D=28
M672 1957 363 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=96880 $Y=55910 $D=28
M673 391 359 1957 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=97200 $Y=55910 $D=28
M674 1958 376 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=101680 $Y=75490 $D=28
M675 372 387 1958 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=102000 $Y=75490 $D=28
M676 1959 438 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=107280 $Y=61090 $D=28
M677 414 833 1959 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=107600 $Y=61090 $D=28
M678 1960 476 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=114080 $Y=63110 $D=28
M679 426 429 1960 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=114400 $Y=63110 $D=28
M680 1961 448 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=114480 $Y=55910 $D=28
M681 838 433 1961 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=114800 $Y=55910 $D=28
M682 1962 443 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=116080 $Y=55910 $D=28
M683 430 838 1962 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=116400 $Y=55910 $D=28
M684 1963 443 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=117680 $Y=63110 $D=28
M685 439 429 1963 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=118000 $Y=63110 $D=28
M686 1964 477 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=121680 $Y=25090 $D=28
M687 427 469 1964 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=122000 $Y=25090 $D=28
M688 1965 456 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=122480 $Y=32290 $D=28
M689 477 471 1965 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=122800 $Y=32290 $D=28
M690 1966 457 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=123280 $Y=55910 $D=28
M691 844 463 1966 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=123600 $Y=55910 $D=28
M692 1967 844 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=126480 $Y=55910 $D=28
M693 481 460 1967 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=126800 $Y=55910 $D=28
M694 1968 502 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=132880 $Y=53890 $D=28
M695 520 524 1968 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=133200 $Y=53890 $D=28
M696 1969 515 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=133680 $Y=32290 $D=28
M697 519 488 1969 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=134000 $Y=32290 $D=28
M698 1970 559 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=138080 $Y=63110 $D=28
M699 560 608 1970 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=138400 $Y=63110 $D=28
M700 1971 558 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=140080 $Y=27110 $D=28
M701 522 853 1971 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=140400 $Y=27110 $D=28
M702 1972 548 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=143680 $Y=68290 $D=28
M703 854 562 1972 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=144000 $Y=68290 $D=28
M704 1973 601 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=147680 $Y=53890 $D=28
M705 557 669 1973 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=148000 $Y=53890 $D=28
M706 1974 602 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=149680 $Y=61090 $D=28
M707 626 595 1974 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=150000 $Y=61090 $D=28
M708 1975 609 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=154480 $Y=61090 $D=28
M709 614 622 1975 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=154800 $Y=61090 $D=28
M710 1976 625 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=157680 $Y=48710 $D=28
M711 624 642 1976 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=158000 $Y=48710 $D=28
M712 1977 632 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=161680 $Y=41510 $D=28
M713 633 639 1977 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=162000 $Y=41510 $D=28
M714 1978 617 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=164480 $Y=68290 $D=28
M715 692 657 1978 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=164800 $Y=68290 $D=28
M716 1979 710 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=166480 $Y=46690 $D=28
M717 712 669 1979 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=166800 $Y=46690 $D=28
M718 1980 576 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=166480 $Y=63110 $D=28
M719 679 670 1980 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=166800 $Y=63110 $D=28
M720 1981 724 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=166880 $Y=41510 $D=28
M721 676 671 1981 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=167200 $Y=41510 $D=28
M722 1982 685 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=167280 $Y=55910 $D=28
M723 713 673 1982 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=167600 $Y=55910 $D=28
M724 1983 726 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=167680 $Y=39490 $D=28
M725 724 675 1983 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=168000 $Y=39490 $D=28
M726 1984 684 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=170080 $Y=63110 $D=28
M727 695 677 1984 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=170400 $Y=63110 $D=28
M728 1985 696 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=171680 $Y=63110 $D=28
M729 785 636 1985 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=172000 $Y=63110 $D=28
M730 1986 732 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=173280 $Y=61090 $D=28
M731 863 707 1986 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=173600 $Y=61090 $D=28
M732 1987 683 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=174480 $Y=34310 $D=28
M733 735 709 1987 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=174800 $Y=34310 $D=28
M734 1988 723 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=175280 $Y=25090 $D=28
M735 715 761 1988 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=175600 $Y=25090 $D=28
M736 1989 652 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=175680 $Y=63110 $D=28
M737 736 744 1989 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=176000 $Y=63110 $D=28
M738 1990 717 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=176880 $Y=25090 $D=28
M739 723 748 1990 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=177200 $Y=25090 $D=28
M740 1991 749 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=179280 $Y=39490 $D=28
M741 752 742 1991 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=179600 $Y=39490 $D=28
M742 1992 759 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=182880 $Y=39490 $D=28
M743 865 778 1992 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=183200 $Y=39490 $D=28
M744 VSS 10 1993 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=10860 $Y=13090 $D=28
M745 798 11 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=11440 $Y=12850 $D=28
M746 VSS 1993 798 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=11920 $Y=12850 $D=28
M747 VSS 25 1995 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=12060 $Y=61090 $D=28
M748 24 23 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=12640 $Y=61090 $D=28
M749 VSS 1995 24 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=13120 $Y=61090 $D=28
M750 VSS 41 1997 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=14060 $Y=61090 $D=28
M751 18 23 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=14640 $Y=61090 $D=28
M752 VSS 1997 18 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=15120 $Y=61090 $D=28
M753 VSS 28 1999 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=14860 $Y=39490 $D=28
M754 801 23 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=15440 $Y=39490 $D=28
M755 VSS 1999 801 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=15920 $Y=39490 $D=28
M756 VSS 122 2001 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=30060 $Y=17890 $D=28
M757 95 11 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=30640 $Y=17890 $D=28
M758 VSS 2001 95 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=31120 $Y=17890 $D=28
M759 VSS 817 2003 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=59660 $Y=17890 $D=28
M760 226 11 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=60240 $Y=17890 $D=28
M761 VSS 2003 226 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=60720 $Y=17890 $D=28
M762 VSS 257 2005 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=69660 $Y=20290 $D=28
M763 261 271 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=70240 $Y=20050 $D=28
M764 VSS 2005 261 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=70720 $Y=20050 $D=28
M765 VSS 217 2007 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=71660 $Y=25090 $D=28
M766 274 148 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=72240 $Y=25090 $D=28
M767 VSS 2007 274 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=72720 $Y=25090 $D=28
M768 VSS 826 2009 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=76860 $Y=20290 $D=28
M769 827 300 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=77440 $Y=20050 $D=28
M770 VSS 2009 827 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=77920 $Y=20050 $D=28
M771 VSS 370 2011 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=104860 $Y=34690 $D=28
M772 386 409 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=105440 $Y=34450 $D=28
M773 VSS 2011 386 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=105920 $Y=34450 $D=28
M774 VSS 573 2013 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=145660 $Y=32290 $D=28
M775 577 582 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=146240 $Y=32290 $D=28
M776 VSS 2013 577 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=146720 $Y=32290 $D=28
M777 VSS 634 2015 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=153660 $Y=49090 $D=28
M778 613 592 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=154240 $Y=48850 $D=28
M779 VSS 2015 613 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=154720 $Y=48850 $D=28
M780 VSS 663 2017 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=156060 $Y=41890 $D=28
M781 647 592 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=156640 $Y=41650 $D=28
M782 VSS 2017 647 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=157120 $Y=41650 $D=28
M783 VSS 865 2019 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55754e-14 as=1.655e-13 pd=6.39692e-07 ps=1.76e-06 nrd=1.14825 nrs=3.41942 sa=3.7e-07 sb=1.3e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=182860 $Y=27490 $D=28
M784 868 681 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.28e-14 as=1.16203e-13 pd=8.2e-07 ps=1.33754e-06 nrd=0.391304 nrs=0.549164 sa=5.79565e-07 sb=7.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=183440 $Y=27250 $D=28
M785 VSS 2019 868 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.19259e-13 as=8.28e-14 pd=1.42259e-06 ps=8.2e-07 nrd=0.563607 nrs=0.391304 sa=1.05957e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=183920 $Y=27250 $D=28
M786 VSS 79 2022 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=25210 $Y=62990 $D=28
M787 2022 79 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=25690 $Y=62990 $D=28
M788 VSS 79 2022 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=26170 $Y=62990 $D=28
M789 2021 110 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=26730 $Y=62830 $D=28
M790 96 2021 2022 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=27920 $Y=62790 $D=28
M791 2022 2021 96 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=28400 $Y=62790 $D=28
M792 96 2021 2022 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=28880 $Y=62790 $D=28
M793 2023 110 96 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=29360 $Y=62790 $D=28
M794 96 110 2023 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=29840 $Y=62790 $D=28
M795 2023 110 96 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=30320 $Y=62790 $D=28
M796 VSS 2022 2023 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=30860 $Y=62790 $D=28
M797 2023 2022 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=31340 $Y=62790 $D=28
M798 VSS 2022 2023 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=31820 $Y=62790 $D=28
M799 VSS 86 2025 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=25210 $Y=68290 $D=28
M800 2025 86 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=25690 $Y=68290 $D=28
M801 VSS 86 2025 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=26170 $Y=68290 $D=28
M802 2024 79 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=26730 $Y=68290 $D=28
M803 73 2024 2025 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=27920 $Y=68510 $D=28
M804 2025 2024 73 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=28400 $Y=68510 $D=28
M805 73 2024 2025 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=28880 $Y=68510 $D=28
M806 2026 79 73 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=29360 $Y=68510 $D=28
M807 73 79 2026 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=29840 $Y=68510 $D=28
M808 2026 79 73 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=30320 $Y=68510 $D=28
M809 VSS 2025 2026 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=30860 $Y=68510 $D=28
M810 2026 2025 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=31340 $Y=68510 $D=28
M811 VSS 2025 2026 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=31820 $Y=68510 $D=28
M812 VSS 141 2028 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=38410 $Y=26990 $D=28
M813 2028 141 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=38890 $Y=26990 $D=28
M814 VSS 141 2028 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=39370 $Y=26990 $D=28
M815 2027 163 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=39930 $Y=26830 $D=28
M816 165 2027 2028 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=41120 $Y=26790 $D=28
M817 2028 2027 165 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=41600 $Y=26790 $D=28
M818 165 2027 2028 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=42080 $Y=26790 $D=28
M819 2029 163 165 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=42560 $Y=26790 $D=28
M820 165 163 2029 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=43040 $Y=26790 $D=28
M821 2029 163 165 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=43520 $Y=26790 $D=28
M822 VSS 2028 2029 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=44060 $Y=26790 $D=28
M823 2029 2028 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=44540 $Y=26790 $D=28
M824 VSS 2028 2029 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=45020 $Y=26790 $D=28
M825 VSS 135 2031 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=39210 $Y=32290 $D=28
M826 2031 135 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=39690 $Y=32290 $D=28
M827 VSS 135 2031 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=40170 $Y=32290 $D=28
M828 2030 123 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=40730 $Y=32290 $D=28
M829 199 2030 2031 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=41920 $Y=32510 $D=28
M830 2031 2030 199 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=42400 $Y=32510 $D=28
M831 199 2030 2031 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=42880 $Y=32510 $D=28
M832 2032 123 199 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=43360 $Y=32510 $D=28
M833 199 123 2032 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=43840 $Y=32510 $D=28
M834 2032 123 199 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=44320 $Y=32510 $D=28
M835 VSS 2031 2032 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=44860 $Y=32510 $D=28
M836 2032 2031 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=45340 $Y=32510 $D=28
M837 VSS 2031 2032 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=45820 $Y=32510 $D=28
M838 VSS 192 2034 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=44810 $Y=34190 $D=28
M839 2034 192 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=45290 $Y=34190 $D=28
M840 VSS 192 2034 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=45770 $Y=34190 $D=28
M841 2033 163 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=46330 $Y=34030 $D=28
M842 144 2033 2034 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=47520 $Y=33990 $D=28
M843 2034 2033 144 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=48000 $Y=33990 $D=28
M844 144 2033 2034 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=48480 $Y=33990 $D=28
M845 2035 163 144 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=48960 $Y=33990 $D=28
M846 144 163 2035 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=49440 $Y=33990 $D=28
M847 2035 163 144 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=49920 $Y=33990 $D=28
M848 VSS 2034 2035 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=50460 $Y=33990 $D=28
M849 2035 2034 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=50940 $Y=33990 $D=28
M850 VSS 2034 2035 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=51420 $Y=33990 $D=28
M851 VSS 49 2037 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=47210 $Y=26990 $D=28
M852 2037 49 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=47690 $Y=26990 $D=28
M853 VSS 49 2037 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=48170 $Y=26990 $D=28
M854 2036 113 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=48730 $Y=26830 $D=28
M855 203 2036 2037 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=49920 $Y=26790 $D=28
M856 2037 2036 203 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=50400 $Y=26790 $D=28
M857 203 2036 2037 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=50880 $Y=26790 $D=28
M858 2038 113 203 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=51360 $Y=26790 $D=28
M859 203 113 2038 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=51840 $Y=26790 $D=28
M860 2038 113 203 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=52320 $Y=26790 $D=28
M861 VSS 2037 2038 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=52860 $Y=26790 $D=28
M862 2038 2037 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=53340 $Y=26790 $D=28
M863 VSS 2037 2038 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=53820 $Y=26790 $D=28
M864 VSS 135 2040 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=55610 $Y=46690 $D=28
M865 2040 135 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=56090 $Y=46690 $D=28
M866 VSS 135 2040 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=56570 $Y=46690 $D=28
M867 2039 123 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=57130 $Y=46690 $D=28
M868 285 2039 2040 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=58320 $Y=46910 $D=28
M869 2040 2039 285 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=58800 $Y=46910 $D=28
M870 285 2039 2040 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=59280 $Y=46910 $D=28
M871 2041 123 285 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=59760 $Y=46910 $D=28
M872 285 123 2041 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=60240 $Y=46910 $D=28
M873 2041 123 285 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=60720 $Y=46910 $D=28
M874 VSS 2040 2041 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=61260 $Y=46910 $D=28
M875 2041 2040 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=61740 $Y=46910 $D=28
M876 VSS 2040 2041 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=62220 $Y=46910 $D=28
M877 VSS 272 2043 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=60010 $Y=75490 $D=28
M878 2043 272 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=60490 $Y=75490 $D=28
M879 VSS 272 2043 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=60970 $Y=75490 $D=28
M880 2042 268 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=61530 $Y=75490 $D=28
M881 819 2042 2043 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=62720 $Y=75710 $D=28
M882 2043 2042 819 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=63200 $Y=75710 $D=28
M883 819 2042 2043 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=63680 $Y=75710 $D=28
M884 2044 268 819 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=64160 $Y=75710 $D=28
M885 819 268 2044 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=64640 $Y=75710 $D=28
M886 2044 268 819 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=65120 $Y=75710 $D=28
M887 VSS 2043 2044 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=65660 $Y=75710 $D=28
M888 2044 2043 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=66140 $Y=75710 $D=28
M889 VSS 2043 2044 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=66620 $Y=75710 $D=28
M890 VSS 289 2046 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=60410 $Y=70190 $D=28
M891 2046 289 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=60890 $Y=70190 $D=28
M892 VSS 289 2046 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=61370 $Y=70190 $D=28
M893 2045 819 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=61930 $Y=70030 $D=28
M894 238 2045 2046 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=63120 $Y=69990 $D=28
M895 2046 2045 238 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=63600 $Y=69990 $D=28
M896 238 2045 2046 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=64080 $Y=69990 $D=28
M897 2047 819 238 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=64560 $Y=69990 $D=28
M898 238 819 2047 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=65040 $Y=69990 $D=28
M899 2047 819 238 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=65520 $Y=69990 $D=28
M900 VSS 2046 2047 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=66060 $Y=69990 $D=28
M901 2047 2046 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=66540 $Y=69990 $D=28
M902 VSS 2046 2047 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=67020 $Y=69990 $D=28
M903 VSS 239 2049 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=65210 $Y=61090 $D=28
M904 2049 239 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=65690 $Y=61090 $D=28
M905 VSS 239 2049 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=66170 $Y=61090 $D=28
M906 2048 248 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=66730 $Y=61090 $D=28
M907 253 2048 2049 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=67920 $Y=61310 $D=28
M908 2049 2048 253 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=68400 $Y=61310 $D=28
M909 253 2048 2049 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=68880 $Y=61310 $D=28
M910 2050 248 253 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=69360 $Y=61310 $D=28
M911 253 248 2050 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=69840 $Y=61310 $D=28
M912 2050 248 253 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=70320 $Y=61310 $D=28
M913 VSS 2049 2050 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=70860 $Y=61310 $D=28
M914 2050 2049 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=71340 $Y=61310 $D=28
M915 VSS 2049 2050 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=71820 $Y=61310 $D=28
M916 VSS 49 2052 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=67210 $Y=26990 $D=28
M917 2052 49 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=67690 $Y=26990 $D=28
M918 VSS 49 2052 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=68170 $Y=26990 $D=28
M919 2051 170 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=68730 $Y=26830 $D=28
M920 212 2051 2052 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=69920 $Y=26790 $D=28
M921 2052 2051 212 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=70400 $Y=26790 $D=28
M922 212 2051 2052 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=70880 $Y=26790 $D=28
M923 2053 170 212 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=71360 $Y=26790 $D=28
M924 212 170 2053 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=71840 $Y=26790 $D=28
M925 2053 170 212 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=72320 $Y=26790 $D=28
M926 VSS 2052 2053 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=72860 $Y=26790 $D=28
M927 2053 2052 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=73340 $Y=26790 $D=28
M928 VSS 2052 2053 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=73820 $Y=26790 $D=28
M929 VSS 254 2055 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=67210 $Y=32290 $D=28
M930 2055 254 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=67690 $Y=32290 $D=28
M931 VSS 254 2055 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=68170 $Y=32290 $D=28
M932 2054 170 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=68730 $Y=32290 $D=28
M933 267 2054 2055 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=69920 $Y=32510 $D=28
M934 2055 2054 267 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=70400 $Y=32510 $D=28
M935 267 2054 2055 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=70880 $Y=32510 $D=28
M936 2056 170 267 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=71360 $Y=32510 $D=28
M937 267 170 2056 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=71840 $Y=32510 $D=28
M938 2056 170 267 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=72320 $Y=32510 $D=28
M939 VSS 2055 2056 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=72860 $Y=32510 $D=28
M940 2056 2055 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=73340 $Y=32510 $D=28
M941 VSS 2055 2056 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=73820 $Y=32510 $D=28
M942 VSS 176 2058 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=79610 $Y=41390 $D=28
M943 2058 176 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=80090 $Y=41390 $D=28
M944 VSS 176 2058 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=80570 $Y=41390 $D=28
M945 2057 307 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=81130 $Y=41230 $D=28
M946 313 2057 2058 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=82320 $Y=41190 $D=28
M947 2058 2057 313 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=82800 $Y=41190 $D=28
M948 313 2057 2058 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=83280 $Y=41190 $D=28
M949 2059 307 313 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=83760 $Y=41190 $D=28
M950 313 307 2059 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=84240 $Y=41190 $D=28
M951 2059 307 313 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=84720 $Y=41190 $D=28
M952 VSS 2058 2059 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=85260 $Y=41190 $D=28
M953 2059 2058 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=85740 $Y=41190 $D=28
M954 VSS 2058 2059 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=86220 $Y=41190 $D=28
M955 VSS 354 2061 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=98010 $Y=41390 $D=28
M956 2061 354 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=98490 $Y=41390 $D=28
M957 VSS 354 2061 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=98970 $Y=41390 $D=28
M958 2060 367 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=99530 $Y=41230 $D=28
M959 419 2060 2061 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-15 $X=100720 $Y=41190 $D=28
M960 2061 2060 419 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-15 $X=101200 $Y=41190 $D=28
M961 419 2060 2061 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=6e-15 $X=101680 $Y=41190 $D=28
M962 2062 367 419 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=6e-15 $X=102160 $Y=41190 $D=28
M963 419 367 2062 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=6e-15 $X=102640 $Y=41190 $D=28
M964 2062 367 419 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=6e-15 $X=103120 $Y=41190 $D=28
M965 VSS 2061 2062 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=103660 $Y=41190 $D=28
M966 2062 2061 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=104140 $Y=41190 $D=28
M967 VSS 2061 2062 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=104620 $Y=41190 $D=28
M968 VSS 909 2064 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=98410 $Y=70190 $D=28
M969 2064 909 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=98890 $Y=70190 $D=28
M970 VSS 909 2064 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=99370 $Y=70190 $D=28
M971 2063 383 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=99930 $Y=70030 $D=28
M972 378 2063 2064 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=101120 $Y=69990 $D=28
M973 2064 2063 378 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=101600 $Y=69990 $D=28
M974 378 2063 2064 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=4e-15 $X=102080 $Y=69990 $D=28
M975 2065 383 378 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-14 $X=102560 $Y=69990 $D=28
M976 378 383 2065 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-14 $X=103040 $Y=69990 $D=28
M977 2065 383 378 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-14 $X=103520 $Y=69990 $D=28
M978 VSS 2064 2065 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-14 $X=104060 $Y=69990 $D=28
M979 2065 2064 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-15 $X=104540 $Y=69990 $D=28
M980 VSS 2064 2065 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-15 $X=105020 $Y=69990 $D=28
M981 VSS 481 2067 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=121210 $Y=61090 $D=28
M982 2067 481 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=121690 $Y=61090 $D=28
M983 VSS 481 2067 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=122170 $Y=61090 $D=28
M984 2066 464 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=7.2e-15 $X=122730 $Y=61090 $D=28
M985 487 2066 2067 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=123920 $Y=61310 $D=28
M986 2067 2066 487 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=124400 $Y=61310 $D=28
M987 487 2066 2067 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=124880 $Y=61310 $D=28
M988 2068 464 487 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=125360 $Y=61310 $D=28
M989 487 464 2068 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=125840 $Y=61310 $D=28
M990 2068 464 487 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=126320 $Y=61310 $D=28
M991 VSS 2067 2068 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=126860 $Y=61310 $D=28
M992 2068 2067 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=127340 $Y=61310 $D=28
M993 VSS 2067 2068 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=127820 $Y=61310 $D=28
M994 VSS 578 2070 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=144810 $Y=62990 $D=28
M995 2070 578 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=145290 $Y=62990 $D=28
M996 VSS 578 2070 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=145770 $Y=62990 $D=28
M997 2069 583 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=146330 $Y=62830 $D=28
M998 590 2069 2070 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=147520 $Y=62790 $D=28
M999 2070 2069 590 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=148000 $Y=62790 $D=28
M1000 590 2069 2070 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=148480 $Y=62790 $D=28
M1001 2071 583 590 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=148960 $Y=62790 $D=28
M1002 590 583 2071 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=149440 $Y=62790 $D=28
M1003 2071 583 590 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=149920 $Y=62790 $D=28
M1004 VSS 2070 2071 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=150460 $Y=62790 $D=28
M1005 2071 2070 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=150940 $Y=62790 $D=28
M1006 VSS 2070 2071 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=151420 $Y=62790 $D=28
M1007 VSS 676 2073 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=168010 $Y=46690 $D=28
M1008 2073 676 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=168490 $Y=46690 $D=28
M1009 VSS 676 2073 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=168970 $Y=46690 $D=28
M1010 2072 702 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=169530 $Y=46690 $D=28
M1011 700 2072 2073 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=170720 $Y=46910 $D=28
M1012 2073 2072 700 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-14 $X=171200 $Y=46910 $D=28
M1013 700 2072 2073 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-14 $X=171680 $Y=46910 $D=28
M1014 2074 702 700 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-14 $X=172160 $Y=46910 $D=28
M1015 700 702 2074 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=172640 $Y=46910 $D=28
M1016 2074 702 700 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=173120 $Y=46910 $D=28
M1017 VSS 2073 2074 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=173660 $Y=46910 $D=28
M1018 2074 2073 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=174140 $Y=46910 $D=28
M1019 VSS 2073 2074 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=174620 $Y=46910 $D=28
M1020 VSS 715 2076 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=181210 $Y=32290 $D=28
M1021 2076 715 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=181690 $Y=32290 $D=28
M1022 VSS 715 2076 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7663e-13 as=1.296e-13 pd=1.24851e-06 ps=1.08e-06 nrd=0.340721 nrs=0.25 sa=1.28e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=182170 $Y=32290 $D=28
M1023 2075 764 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.696e-13 as=2.15881e-13 pd=2.4e-06 ps=1.52596e-06 nrd=0.34814 nrs=0.278772 sa=1.57091e-06 sb=3.06364e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=182730 $Y=32290 $D=28
M1024 743 2075 2076 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.084e-13 pd=1.06e-06 ps=2.04e-06 nrd=0.257143 nrs=0.425306 sa=2.97714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=183920 $Y=32510 $D=28
M1025 2076 2075 743 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.77714e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=184400 $Y=32510 $D=28
M1026 743 2075 2076 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.25771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=184880 $Y=32510 $D=28
M1027 2077 764 743 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.73771e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=185360 $Y=32510 $D=28
M1028 743 764 2077 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=185840 $Y=32510 $D=28
M1029 2077 764 743 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47e-13 as=1.26e-13 pd=1.12e-06 ps=1.06e-06 nrd=0.3 nrs=0.257143 sa=2e-06 sb=1.82e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=186320 $Y=32510 $D=28
M1030 VSS 2076 2077 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.47e-13 pd=1.06e-06 ps=1.12e-06 nrd=0.257143 nrs=0.3 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=186860 $Y=32510 $D=28
M1031 2077 2076 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=187340 $Y=32510 $D=28
M1032 VSS 2076 2077 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.24e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.457143 nrs=0.257143 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=187820 $Y=32510 $D=28
M1033 2079 52 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=18940 $Y=32290 $D=28
M1034 VSS 52 2079 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=19420 $Y=32290 $D=28
M1035 2079 52 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=19900 $Y=32290 $D=28
M1036 VSS 52 2079 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=20380 $Y=32290 $D=28
M1037 2078 70 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=20940 $Y=32290 $D=28
M1038 26 70 2079 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=21900 $Y=32410 $D=28
M1039 2079 70 26 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=22380 $Y=32410 $D=28
M1040 26 70 2079 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=22860 $Y=32410 $D=28
M1041 2080 2078 26 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=23340 $Y=32410 $D=28
M1042 26 2078 2080 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=23820 $Y=32410 $D=28
M1043 2080 2078 26 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=24300 $Y=32410 $D=28
M1044 VSS 2079 2080 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=24780 $Y=32410 $D=28
M1045 2080 2079 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=25260 $Y=32410 $D=28
M1046 VSS 2079 2080 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=25740 $Y=32410 $D=28
M1047 2082 109 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=25340 $Y=53890 $D=28
M1048 VSS 109 2082 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=25820 $Y=53890 $D=28
M1049 2082 109 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=26300 $Y=53890 $D=28
M1050 VSS 109 2082 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=26780 $Y=53890 $D=28
M1051 2081 99 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=27340 $Y=53890 $D=28
M1052 92 99 2082 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=28300 $Y=54010 $D=28
M1053 2082 99 92 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=28780 $Y=54010 $D=28
M1054 92 99 2082 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=29260 $Y=54010 $D=28
M1055 2083 2081 92 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=29740 $Y=54010 $D=28
M1056 92 2081 2083 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=30220 $Y=54010 $D=28
M1057 2083 2081 92 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=30700 $Y=54010 $D=28
M1058 VSS 2082 2083 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=31180 $Y=54010 $D=28
M1059 2083 2082 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=31660 $Y=54010 $D=28
M1060 VSS 2082 2083 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=32140 $Y=54010 $D=28
M1061 2085 211 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=31740 $Y=55960 $D=28
M1062 VSS 211 2085 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=32220 $Y=55960 $D=28
M1063 2085 211 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=32700 $Y=55960 $D=28
M1064 VSS 211 2085 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=33180 $Y=55960 $D=28
M1065 2084 160 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=33740 $Y=55630 $D=28
M1066 99 160 2085 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=34700 $Y=55670 $D=28
M1067 2085 160 99 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=35180 $Y=55670 $D=28
M1068 99 160 2085 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=35660 $Y=55670 $D=28
M1069 2086 2084 99 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=36140 $Y=55670 $D=28
M1070 99 2084 2086 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=36620 $Y=55670 $D=28
M1071 2086 2084 99 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=37100 $Y=55670 $D=28
M1072 VSS 2085 2086 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=37580 $Y=55670 $D=28
M1073 2086 2085 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=38060 $Y=55670 $D=28
M1074 VSS 2085 2086 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=38540 $Y=55670 $D=28
M1075 2088 140 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=46540 $Y=19960 $D=28
M1076 VSS 140 2088 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=47020 $Y=19960 $D=28
M1077 2088 140 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=47500 $Y=19960 $D=28
M1078 VSS 140 2088 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=47980 $Y=19960 $D=28
M1079 2087 173 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=48540 $Y=19630 $D=28
M1080 188 173 2088 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=49500 $Y=19670 $D=28
M1081 2088 173 188 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=49980 $Y=19670 $D=28
M1082 188 173 2088 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=50460 $Y=19670 $D=28
M1083 2089 2087 188 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=50940 $Y=19670 $D=28
M1084 188 2087 2089 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=51420 $Y=19670 $D=28
M1085 2089 2087 188 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=51900 $Y=19670 $D=28
M1086 VSS 2088 2089 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=52380 $Y=19670 $D=28
M1087 2089 2088 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=52860 $Y=19670 $D=28
M1088 VSS 2088 2089 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=53340 $Y=19670 $D=28
M1089 2091 201 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=52940 $Y=48760 $D=28
M1090 VSS 201 2091 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=53420 $Y=48760 $D=28
M1091 2091 201 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=53900 $Y=48760 $D=28
M1092 VSS 201 2091 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=54380 $Y=48760 $D=28
M1093 2090 195 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=54940 $Y=48430 $D=28
M1094 213 195 2091 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=55900 $Y=48470 $D=28
M1095 2091 195 213 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=56380 $Y=48470 $D=28
M1096 213 195 2091 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=56860 $Y=48470 $D=28
M1097 2092 2090 213 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=57340 $Y=48470 $D=28
M1098 213 2090 2092 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=57820 $Y=48470 $D=28
M1099 2092 2090 213 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=58300 $Y=48470 $D=28
M1100 VSS 2091 2092 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=58780 $Y=48470 $D=28
M1101 2092 2091 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=59260 $Y=48470 $D=28
M1102 VSS 2091 2092 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=59740 $Y=48470 $D=28
M1103 2094 210 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=54140 $Y=61090 $D=28
M1104 VSS 210 2094 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=54620 $Y=61090 $D=28
M1105 2094 210 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=55100 $Y=61090 $D=28
M1106 VSS 210 2094 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=55580 $Y=61090 $D=28
M1107 2093 220 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=56140 $Y=61090 $D=28
M1108 230 220 2094 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=57100 $Y=61210 $D=28
M1109 2094 220 230 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=57580 $Y=61210 $D=28
M1110 230 220 2094 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=58060 $Y=61210 $D=28
M1111 2095 2093 230 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=58540 $Y=61210 $D=28
M1112 230 2093 2095 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=59020 $Y=61210 $D=28
M1113 2095 2093 230 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=59500 $Y=61210 $D=28
M1114 VSS 2094 2095 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=59980 $Y=61210 $D=28
M1115 2095 2094 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=60460 $Y=61210 $D=28
M1116 VSS 2094 2095 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=60940 $Y=61210 $D=28
M1117 2097 135 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=59340 $Y=27160 $D=28
M1118 VSS 135 2097 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=59820 $Y=27160 $D=28
M1119 2097 135 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=60300 $Y=27160 $D=28
M1120 VSS 135 2097 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=60780 $Y=27160 $D=28
M1121 2096 231 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=61340 $Y=26830 $D=28
M1122 236 231 2097 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=62300 $Y=26870 $D=28
M1123 2097 231 236 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=62780 $Y=26870 $D=28
M1124 236 231 2097 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=63260 $Y=26870 $D=28
M1125 2098 2096 236 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=63740 $Y=26870 $D=28
M1126 236 2096 2098 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=64220 $Y=26870 $D=28
M1127 2098 2096 236 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=64700 $Y=26870 $D=28
M1128 VSS 2097 2098 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=65180 $Y=26870 $D=28
M1129 2098 2097 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=65660 $Y=26870 $D=28
M1130 VSS 2097 2098 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=66140 $Y=26870 $D=28
M1131 2100 263 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=60140 $Y=39490 $D=28
M1132 VSS 263 2100 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=60620 $Y=39490 $D=28
M1133 2100 263 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=61100 $Y=39490 $D=28
M1134 VSS 263 2100 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=61580 $Y=39490 $D=28
M1135 2099 228 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=62140 $Y=39490 $D=28
M1136 237 228 2100 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=63100 $Y=39610 $D=28
M1137 2100 228 237 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=63580 $Y=39610 $D=28
M1138 237 228 2100 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=64060 $Y=39610 $D=28
M1139 2101 2099 237 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=64540 $Y=39610 $D=28
M1140 237 2099 2101 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=65020 $Y=39610 $D=28
M1141 2101 2099 237 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=65500 $Y=39610 $D=28
M1142 VSS 2100 2101 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=65980 $Y=39610 $D=28
M1143 2101 2100 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=66460 $Y=39610 $D=28
M1144 VSS 2100 2101 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=66940 $Y=39610 $D=28
M1145 2103 359 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=86940 $Y=55960 $D=28
M1146 VSS 359 2103 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=87420 $Y=55960 $D=28
M1147 2103 359 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=87900 $Y=55960 $D=28
M1148 VSS 359 2103 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=88380 $Y=55960 $D=28
M1149 2102 352 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=88940 $Y=55630 $D=28
M1150 355 352 2103 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=89900 $Y=55670 $D=28
M1151 2103 352 355 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=90380 $Y=55670 $D=28
M1152 355 352 2103 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=90860 $Y=55670 $D=28
M1153 2104 2102 355 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=91340 $Y=55670 $D=28
M1154 355 2102 2104 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=91820 $Y=55670 $D=28
M1155 2104 2102 355 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=92300 $Y=55670 $D=28
M1156 VSS 2103 2104 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=92780 $Y=55670 $D=28
M1157 2104 2103 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=93260 $Y=55670 $D=28
M1158 VSS 2103 2104 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=93740 $Y=55670 $D=28
M1159 2106 363 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=90940 $Y=53890 $D=28
M1160 VSS 363 2106 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=91420 $Y=53890 $D=28
M1161 2106 363 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=91900 $Y=53890 $D=28
M1162 VSS 363 2106 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=92380 $Y=53890 $D=28
M1163 2105 348 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=92940 $Y=53890 $D=28
M1164 352 348 2106 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=93900 $Y=54010 $D=28
M1165 2106 348 352 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=94380 $Y=54010 $D=28
M1166 352 348 2106 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=94860 $Y=54010 $D=28
M1167 2107 2105 352 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=95340 $Y=54010 $D=28
M1168 352 2105 2107 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=95820 $Y=54010 $D=28
M1169 2107 2105 352 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=96300 $Y=54010 $D=28
M1170 VSS 2106 2107 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=96780 $Y=54010 $D=28
M1171 2107 2106 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=97260 $Y=54010 $D=28
M1172 VSS 2106 2107 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=97740 $Y=54010 $D=28
M1173 2109 398 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=99340 $Y=53890 $D=28
M1174 VSS 398 2109 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=99820 $Y=53890 $D=28
M1175 2109 398 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=100300 $Y=53890 $D=28
M1176 VSS 398 2109 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=100780 $Y=53890 $D=28
M1177 2108 395 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=101340 $Y=53890 $D=28
M1178 380 395 2109 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=102300 $Y=54010 $D=28
M1179 2109 395 380 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=102780 $Y=54010 $D=28
M1180 380 395 2109 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=103260 $Y=54010 $D=28
M1181 2110 2108 380 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=103740 $Y=54010 $D=28
M1182 380 2108 2110 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=104220 $Y=54010 $D=28
M1183 2110 2108 380 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=104700 $Y=54010 $D=28
M1184 VSS 2109 2110 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=105180 $Y=54010 $D=28
M1185 2110 2109 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=105660 $Y=54010 $D=28
M1186 VSS 2109 2110 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=106140 $Y=54010 $D=28
M1187 2112 426 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=108940 $Y=61090 $D=28
M1188 VSS 426 2112 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=109420 $Y=61090 $D=28
M1189 2112 426 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=109900 $Y=61090 $D=28
M1190 VSS 426 2112 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=110380 $Y=61090 $D=28
M1191 2111 415 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=110940 $Y=61090 $D=28
M1192 394 415 2112 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=111900 $Y=61210 $D=28
M1193 2112 415 394 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=112380 $Y=61210 $D=28
M1194 394 415 2112 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=112860 $Y=61210 $D=28
M1195 2113 2111 394 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=113340 $Y=61210 $D=28
M1196 394 2111 2113 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=113820 $Y=61210 $D=28
M1197 2113 2111 394 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=114300 $Y=61210 $D=28
M1198 VSS 2112 2113 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=114780 $Y=61210 $D=28
M1199 2113 2112 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=115260 $Y=61210 $D=28
M1200 VSS 2112 2113 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=115740 $Y=61210 $D=28
M1201 2115 507 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=125340 $Y=25090 $D=28
M1202 VSS 507 2115 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=125820 $Y=25090 $D=28
M1203 2115 507 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=126300 $Y=25090 $D=28
M1204 VSS 507 2115 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=126780 $Y=25090 $D=28
M1205 2114 483 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=127340 $Y=25090 $D=28
M1206 514 483 2115 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=128300 $Y=25210 $D=28
M1207 2115 483 514 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=128780 $Y=25210 $D=28
M1208 514 483 2115 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=129260 $Y=25210 $D=28
M1209 2116 2114 514 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=129740 $Y=25210 $D=28
M1210 514 2114 2116 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=130220 $Y=25210 $D=28
M1211 2116 2114 514 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=130700 $Y=25210 $D=28
M1212 VSS 2115 2116 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=131180 $Y=25210 $D=28
M1213 2116 2115 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=131660 $Y=25210 $D=28
M1214 VSS 2115 2116 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=132140 $Y=25210 $D=28
M1215 2118 498 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=128940 $Y=61090 $D=28
M1216 VSS 498 2118 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=129420 $Y=61090 $D=28
M1217 2118 498 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=129900 $Y=61090 $D=28
M1218 VSS 498 2118 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=130380 $Y=61090 $D=28
M1219 2117 511 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=130940 $Y=61090 $D=28
M1220 521 511 2118 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=131900 $Y=61210 $D=28
M1221 2118 511 521 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=132380 $Y=61210 $D=28
M1222 521 511 2118 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=132860 $Y=61210 $D=28
M1223 2119 2117 521 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=133340 $Y=61210 $D=28
M1224 521 2117 2119 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=133820 $Y=61210 $D=28
M1225 2119 2117 521 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=134300 $Y=61210 $D=28
M1226 VSS 2118 2119 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=134780 $Y=61210 $D=28
M1227 2119 2118 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=135260 $Y=61210 $D=28
M1228 VSS 2118 2119 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=135740 $Y=61210 $D=28
M1229 2121 555 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=137340 $Y=34360 $D=28
M1230 VSS 555 2121 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=137820 $Y=34360 $D=28
M1231 2121 555 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=138300 $Y=34360 $D=28
M1232 VSS 555 2121 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=138780 $Y=34360 $D=28
M1233 2120 542 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=139340 $Y=34030 $D=28
M1234 535 542 2121 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=140300 $Y=34070 $D=28
M1235 2121 542 535 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=140780 $Y=34070 $D=28
M1236 535 542 2121 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=141260 $Y=34070 $D=28
M1237 2122 2120 535 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=141740 $Y=34070 $D=28
M1238 535 2120 2122 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=142220 $Y=34070 $D=28
M1239 2122 2120 535 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=142700 $Y=34070 $D=28
M1240 VSS 2121 2122 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=143180 $Y=34070 $D=28
M1241 2122 2121 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=143660 $Y=34070 $D=28
M1242 VSS 2121 2122 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=144140 $Y=34070 $D=28
M1243 2124 672 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=156140 $Y=70360 $D=28
M1244 VSS 672 2124 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=156620 $Y=70360 $D=28
M1245 2124 672 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=157100 $Y=70360 $D=28
M1246 VSS 672 2124 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=157580 $Y=70360 $D=28
M1247 2123 857 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=158140 $Y=70030 $D=28
M1248 644 857 2124 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=159100 $Y=70070 $D=28
M1249 2124 857 644 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=159580 $Y=70070 $D=28
M1250 644 857 2124 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=160060 $Y=70070 $D=28
M1251 2125 2123 644 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=160540 $Y=70070 $D=28
M1252 644 2123 2125 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=161020 $Y=70070 $D=28
M1253 2125 2123 644 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=161500 $Y=70070 $D=28
M1254 VSS 2124 2125 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=161980 $Y=70070 $D=28
M1255 2125 2124 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=162460 $Y=70070 $D=28
M1256 VSS 2124 2125 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=162940 $Y=70070 $D=28
M1257 2127 861 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=169340 $Y=75490 $D=28
M1258 VSS 861 2127 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=169820 $Y=75490 $D=28
M1259 2127 861 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=170300 $Y=75490 $D=28
M1260 VSS 861 2127 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=170780 $Y=75490 $D=28
M1261 2126 763 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=171340 $Y=75490 $D=28
M1262 705 763 2127 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=172300 $Y=75610 $D=28
M1263 2127 763 705 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=172780 $Y=75610 $D=28
M1264 705 763 2127 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=173260 $Y=75610 $D=28
M1265 2128 2126 705 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=173740 $Y=75610 $D=28
M1266 705 2126 2128 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=174220 $Y=75610 $D=28
M1267 2128 2126 705 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=174700 $Y=75610 $D=28
M1268 VSS 2127 2128 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=175180 $Y=75610 $D=28
M1269 2128 2127 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=175660 $Y=75610 $D=28
M1270 VSS 2127 2128 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=176140 $Y=75610 $D=28
M1271 2130 774 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=179740 $Y=19960 $D=28
M1272 VSS 774 2130 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=180220 $Y=19960 $D=28
M1273 2130 774 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=180700 $Y=19960 $D=28
M1274 VSS 774 2130 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=181180 $Y=19960 $D=28
M1275 2129 787 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=181740 $Y=19630 $D=28
M1276 767 787 2130 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=182700 $Y=19670 $D=28
M1277 2130 787 767 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=183180 $Y=19670 $D=28
M1278 767 787 2130 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=183660 $Y=19670 $D=28
M1279 2131 2129 767 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=184140 $Y=19670 $D=28
M1280 767 2129 2131 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=184620 $Y=19670 $D=28
M1281 2131 2129 767 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=185100 $Y=19670 $D=28
M1282 VSS 2130 2131 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=185580 $Y=19670 $D=28
M1283 2131 2130 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=186060 $Y=19670 $D=28
M1284 VSS 2130 2131 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=186540 $Y=19670 $D=28
M1285 2133 753 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=180940 $Y=55960 $D=28
M1286 VSS 753 2133 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=181420 $Y=55960 $D=28
M1287 2133 753 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=181900 $Y=55960 $D=28
M1288 VSS 753 2133 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=182380 $Y=55960 $D=28
M1289 2132 866 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=182940 $Y=55630 $D=28
M1290 768 866 2133 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=183900 $Y=55670 $D=28
M1291 2133 866 768 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=184380 $Y=55670 $D=28
M1292 768 866 2133 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=184860 $Y=55670 $D=28
M1293 2134 2132 768 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=185340 $Y=55670 $D=28
M1294 768 2132 2134 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=185820 $Y=55670 $D=28
M1295 2134 2132 768 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=186300 $Y=55670 $D=28
M1296 VSS 2133 2134 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=186780 $Y=55670 $D=28
M1297 2134 2133 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=187260 $Y=55670 $D=28
M1298 VSS 2133 2134 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=187740 $Y=55670 $D=28
M1299 2136 738 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=2.49952e-13 pd=9.1e-07 ps=2.05422e-06 nrd=0.327273 nrs=0.826287 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=180940 $Y=63160 $D=28
M1300 VSS 738 2136 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8.4e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=181420 $Y=63160 $D=28
M1301 2136 738 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.32e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=181900 $Y=63160 $D=28
M1302 VSS 738 2136 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43965e-13 as=9.9e-14 pd=1.04854e-06 ps=9.1e-07 nrd=0.475917 nrs=0.327273 sa=1.8e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=182380 $Y=63160 $D=28
M1303 2135 751 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.30344e-13 pd=2.4e-06 ps=1.67766e-06 nrd=0.363636 nrs=0.297448 sa=1.385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.16e-14 panw10=0 $X=182940 $Y=62830 $D=28
M1304 777 751 2136 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=2.304e-13 pd=1.08e-06 ps=2.08e-06 nrd=0.25 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=183900 $Y=62870 $D=28
M1305 2136 751 777 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=184380 $Y=62870 $D=28
M1306 777 751 2136 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=184860 $Y=62870 $D=28
M1307 2137 2135 777 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=1.76e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=185340 $Y=62870 $D=28
M1308 777 2135 2137 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=185820 $Y=62870 $D=28
M1309 2137 2135 777 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=186300 $Y=62870 $D=28
M1310 VSS 2136 2137 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=186780 $Y=62870 $D=28
M1311 2137 2136 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.296e-13 as=1.296e-13 pd=1.08e-06 ps=1.08e-06 nrd=0.25 nrs=0.25 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=187260 $Y=62870 $D=28
M1312 VSS 2136 2137 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.296e-13 pd=2.08e-06 ps=1.08e-06 nrd=0.444444 nrs=0.25 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=187740 $Y=62870 $D=28
M1313 2138 62 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=13960 $Y=27070 $D=28
M1314 33 27 2138 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=14280 $Y=27070 $D=28
M1315 2139 27 33 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=14760 $Y=27070 $D=28
M1316 VSS 62 2139 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=15080 $Y=27070 $D=28
M1317 2140 133 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=15560 $Y=19870 $D=28
M1318 40 39 2140 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=15880 $Y=19870 $D=28
M1319 2141 39 40 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=16360 $Y=19870 $D=28
M1320 VSS 133 2141 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=16680 $Y=19870 $D=28
M1321 2142 65 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=21160 $Y=70270 $D=28
M1322 105 803 2142 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=21480 $Y=70270 $D=28
M1323 2143 803 105 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=21960 $Y=70270 $D=28
M1324 VSS 65 2143 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=22280 $Y=70270 $D=28
M1325 2144 121 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=23160 $Y=68330 $D=28
M1326 85 69 2144 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=23480 $Y=68330 $D=28
M1327 2145 69 85 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=23960 $Y=68330 $D=28
M1328 VSS 121 2145 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=24280 $Y=68330 $D=28
M1329 2146 87 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=25960 $Y=39530 $D=28
M1330 108 145 2146 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=26280 $Y=39530 $D=28
M1331 2147 145 108 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=26760 $Y=39530 $D=28
M1332 VSS 87 2147 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=27080 $Y=39530 $D=28
M1333 2148 138 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=32360 $Y=61130 $D=28
M1334 807 109 2148 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=32680 $Y=61130 $D=28
M1335 2149 109 807 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=33160 $Y=61130 $D=28
M1336 VSS 138 2149 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=33480 $Y=61130 $D=28
M1337 2150 138 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=33160 $Y=68330 $D=28
M1338 890 139 2150 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=33480 $Y=68330 $D=28
M1339 2151 139 890 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=33960 $Y=68330 $D=28
M1340 VSS 138 2151 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=34280 $Y=68330 $D=28
M1341 2152 191 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=34760 $Y=70270 $D=28
M1342 91 238 2152 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=35080 $Y=70270 $D=28
M1343 2153 238 91 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=35560 $Y=70270 $D=28
M1344 VSS 191 2153 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=35880 $Y=70270 $D=28
M1345 2154 125 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=35960 $Y=19870 $D=28
M1346 132 130 2154 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=36280 $Y=19870 $D=28
M1347 2155 130 132 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=36760 $Y=19870 $D=28
M1348 VSS 125 2155 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=37080 $Y=19870 $D=28
M1349 2156 109 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=39160 $Y=63070 $D=28
M1350 161 139 2156 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=39480 $Y=63070 $D=28
M1351 2157 139 161 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=39960 $Y=63070 $D=28
M1352 VSS 109 2157 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=40280 $Y=63070 $D=28
M1353 2158 205 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=55960 $Y=19870 $D=28
M1354 815 167 2158 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=56280 $Y=19870 $D=28
M1355 2159 167 815 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=56760 $Y=19870 $D=28
M1356 VSS 205 2159 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=57080 $Y=19870 $D=28
M1357 2160 818 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=61960 $Y=61130 $D=28
M1358 233 230 2160 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=62280 $Y=61130 $D=28
M1359 2161 230 233 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=62760 $Y=61130 $D=28
M1360 VSS 818 2161 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=63080 $Y=61130 $D=28
M1361 2162 821 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=68360 $Y=70270 $D=28
M1362 904 823 2162 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=68680 $Y=70270 $D=28
M1363 2163 823 904 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=69160 $Y=70270 $D=28
M1364 VSS 821 2163 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=69480 $Y=70270 $D=28
M1365 2164 342 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=90360 $Y=75530 $D=28
M1366 361 323 2164 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=90680 $Y=75530 $D=28
M1367 2165 323 361 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=91160 $Y=75530 $D=28
M1368 VSS 342 2165 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=91480 $Y=75530 $D=28
M1369 2166 360 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=98360 $Y=55870 $D=28
M1370 375 363 2166 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=98680 $Y=55870 $D=28
M1371 2167 363 375 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=99160 $Y=55870 $D=28
M1372 VSS 360 2167 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=99480 $Y=55870 $D=28
M1373 2168 360 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=100760 $Y=61130 $D=28
M1374 379 359 2168 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=101080 $Y=61130 $D=28
M1375 2169 359 379 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=101560 $Y=61130 $D=28
M1376 VSS 360 2169 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=101880 $Y=61130 $D=28
M1377 2170 448 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=115560 $Y=63070 $D=28
M1378 432 433 2170 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=115880 $Y=63070 $D=28
M1379 2171 433 432 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=116360 $Y=63070 $D=28
M1380 VSS 448 2171 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=116680 $Y=63070 $D=28
M1381 2172 450 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=117560 $Y=32330 $D=28
M1382 445 441 2172 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=117880 $Y=32330 $D=28
M1383 2173 441 445 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=118360 $Y=32330 $D=28
M1384 VSS 450 2173 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=118680 $Y=32330 $D=28
M1385 2174 845 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=127160 $Y=41470 $D=28
M1386 502 480 2174 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=127480 $Y=41470 $D=28
M1387 2175 480 502 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=127960 $Y=41470 $D=28
M1388 VSS 845 2175 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=128280 $Y=41470 $D=28
M1389 2176 493 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=129160 $Y=41470 $D=28
M1390 517 470 2176 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=129480 $Y=41470 $D=28
M1391 2177 470 517 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=129960 $Y=41470 $D=28
M1392 VSS 493 2177 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=130280 $Y=41470 $D=28
M1393 2178 510 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=137160 $Y=46730 $D=28
M1394 512 525 2178 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=137480 $Y=46730 $D=28
M1395 2179 525 512 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=137960 $Y=46730 $D=28
M1396 VSS 510 2179 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=138280 $Y=46730 $D=28
M1397 2180 577 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=145160 $Y=34270 $D=28
M1398 585 571 2180 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=145480 $Y=34270 $D=28
M1399 2181 571 585 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=145960 $Y=34270 $D=28
M1400 VSS 577 2181 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=146280 $Y=34270 $D=28
M1401 2182 613 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=147960 $Y=48670 $D=28
M1402 580 587 2182 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=148280 $Y=48670 $D=28
M1403 2183 587 580 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=148760 $Y=48670 $D=28
M1404 VSS 613 2183 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=149080 $Y=48670 $D=28
M1405 2184 647 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=161160 $Y=48670 $D=28
M1406 649 637 2184 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=161480 $Y=48670 $D=28
M1407 2185 637 649 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=161960 $Y=48670 $D=28
M1408 VSS 647 2185 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=162280 $Y=48670 $D=28
M1409 2186 781 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.95843e-13 pd=8e-07 ps=2.04944e-06 nrd=0.166667 nrs=0.544007 sa=2.7e-07 sb=1.42e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=180760 $Y=39530 $D=28
M1410 779 752 2186 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=6e-14 pd=9.6e-07 ps=8e-07 nrd=0.3 nrs=0.166667 sa=5.9e-07 sb=1.1e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=181080 $Y=39530 $D=28
M1411 2187 752 779 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.08e-13 pd=8e-07 ps=9.6e-07 nrd=0.166667 nrs=0.3 sa=1.07e-06 sb=6.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=181560 $Y=39530 $D=28
M1412 VSS 781 2187 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.14636e-13 as=6e-14 pd=2.05909e-06 ps=8e-07 nrd=0.596212 nrs=0.166667 sa=1.39e-06 sb=3e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=181880 $Y=39530 $D=28
M1413 51 80 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=20920 $Y=63250 $D=28
M1414 2188 51 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=19280 $Y=63110 $D=28
M1415 54 50 2188 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=19600 $Y=63110 $D=28
M1416 847 504 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=129720 $Y=27250 $D=28
M1417 2189 474 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=128080 $Y=27110 $D=28
M1418 504 486 2189 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=128400 $Y=27110 $D=28
M1419 851 527 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=134520 $Y=27250 $D=28
M1420 2190 501 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=132880 $Y=27110 $D=28
M1421 509 469 2190 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=133200 $Y=27110 $D=28
M1422 853 528 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=138920 $Y=27250 $D=28
M1423 2191 505 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=137280 $Y=27110 $D=28
M1424 536 529 2191 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=137600 $Y=27110 $D=28
M1425 569 632 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=146520 $Y=27250 $D=28
M1426 2192 568 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=144880 $Y=27110 $D=28
M1427 554 569 2192 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=145200 $Y=27110 $D=28
M1428 595 581 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=148520 $Y=61090 $D=28
M1429 2193 607 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=146880 $Y=61090 $D=28
M1430 578 595 2193 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=147200 $Y=61090 $D=28
M1431 588 609 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=151720 $Y=56050 $D=28
M1432 2194 597 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=150080 $Y=55910 $D=28
M1433 607 588 2194 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=150400 $Y=55910 $D=28
M1434 629 660 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=163320 $Y=46690 $D=28
M1435 2195 646 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=161680 $Y=46690 $D=28
M1436 660 630 2195 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=162000 $Y=46690 $D=28
M1437 744 746 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.518e-13 pd=1.56e-06 ps=1.58e-06 nrd=0.695652 nrs=0.717391 sa=3.3e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=181720 $Y=53890 $D=28
M1438 2196 746 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.34e-13 pd=8e-07 ps=1.98e-06 nrd=0.166667 nrs=0.65 sa=3.9e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=180080 $Y=53890 $D=28
M1439 734 750 2196 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=7.1e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=180400 $Y=53890 $D=28
M1440 2198 26 2197 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=1.728e-13 pd=7.4e-07 ps=1.72e-06 nrd=0.185185 nrs=0.592593 sa=3.2e-07 sb=1.6437e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=11090 $Y=27120 $D=28
M1441 VSS 47 2198 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21728e-13 as=5.4e-14 pd=1.23972e-06 ps=7.4e-07 nrd=0.417449 nrs=0.185185 sa=6.4e-07 sb=1.54389e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=11410 $Y=27120 $D=28
M1442 2199 33 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.35254e-13 pd=8e-07 ps=1.37746e-06 nrd=0.166667 nrs=0.375704 sa=8.48167e-07 sb=1.288e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=11900 $Y=26930 $D=28
M1443 66 2197 2199 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.104e-13 as=6e-14 pd=1.08e-06 ps=8e-07 nrd=0.306667 nrs=0.166667 sa=1.16817e-06 sb=9.68e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=12220 $Y=26930 $D=28
M1444 2200 2197 66 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.104e-13 pd=8e-07 ps=1.08e-06 nrd=0.166667 nrs=0.306667 sa=1.48017e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=12700 $Y=27050 $D=28
M1445 VSS 33 2200 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.48455e-13 as=6e-14 pd=2.03182e-06 ps=8e-07 nrd=0.690152 nrs=0.166667 sa=1.62933e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=13020 $Y=27050 $D=28
M1446 2202 151 2201 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=1.728e-13 pd=7.4e-07 ps=1.72e-06 nrd=0.185185 nrs=0.592593 sa=3.2e-07 sb=1.6437e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=51090 $Y=61140 $D=28
M1447 VSS 189 2202 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21728e-13 as=5.4e-14 pd=1.23972e-06 ps=7.4e-07 nrd=0.417449 nrs=0.185185 sa=6.4e-07 sb=1.54389e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=51410 $Y=61140 $D=28
M1448 2203 193 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.35254e-13 pd=8e-07 ps=1.37746e-06 nrd=0.166667 nrs=0.375704 sa=8.48167e-07 sb=1.288e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=51900 $Y=61270 $D=28
M1449 340 2201 2203 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.104e-13 as=6e-14 pd=1.08e-06 ps=8e-07 nrd=0.306667 nrs=0.166667 sa=1.16817e-06 sb=9.68e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=52220 $Y=61270 $D=28
M1450 2204 2201 340 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.104e-13 pd=8e-07 ps=1.08e-06 nrd=0.166667 nrs=0.306667 sa=1.48017e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=52700 $Y=61150 $D=28
M1451 VSS 193 2204 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.48455e-13 as=6e-14 pd=2.03182e-06 ps=8e-07 nrd=0.690152 nrs=0.166667 sa=1.62933e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=53020 $Y=61150 $D=28
M1452 2206 215 2205 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=1.728e-13 pd=7.4e-07 ps=1.72e-06 nrd=0.185185 nrs=0.592593 sa=3.2e-07 sb=1.6437e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=62690 $Y=55920 $D=28
M1453 VSS 220 2206 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21728e-13 as=5.4e-14 pd=1.23972e-06 ps=7.4e-07 nrd=0.417449 nrs=0.185185 sa=6.4e-07 sb=1.54389e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=63010 $Y=55920 $D=28
M1454 2207 229 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.35254e-13 pd=8e-07 ps=1.37746e-06 nrd=0.166667 nrs=0.375704 sa=8.48167e-07 sb=1.288e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=63500 $Y=55730 $D=28
M1455 275 2205 2207 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.104e-13 as=6e-14 pd=1.08e-06 ps=8e-07 nrd=0.306667 nrs=0.166667 sa=1.16817e-06 sb=9.68e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=63820 $Y=55730 $D=28
M1456 2208 2205 275 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.104e-13 pd=8e-07 ps=1.08e-06 nrd=0.166667 nrs=0.306667 sa=1.48017e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=64300 $Y=55850 $D=28
M1457 VSS 229 2208 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.48455e-13 as=6e-14 pd=2.03182e-06 ps=8e-07 nrd=0.690152 nrs=0.166667 sa=1.62933e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=64620 $Y=55850 $D=28
M1458 2210 268 2209 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=1.728e-13 pd=7.4e-07 ps=1.72e-06 nrd=0.185185 nrs=0.592593 sa=3.2e-07 sb=1.6437e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=71890 $Y=75540 $D=28
M1459 VSS 272 2210 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21728e-13 as=5.4e-14 pd=1.23972e-06 ps=7.4e-07 nrd=0.417449 nrs=0.185185 sa=6.4e-07 sb=1.54389e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=72210 $Y=75540 $D=28
M1460 2211 277 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.35254e-13 pd=8e-07 ps=1.37746e-06 nrd=0.166667 nrs=0.375704 sa=8.48167e-07 sb=1.288e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=72700 $Y=75670 $D=28
M1461 308 2209 2211 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.104e-13 as=6e-14 pd=1.08e-06 ps=8e-07 nrd=0.306667 nrs=0.166667 sa=1.16817e-06 sb=9.68e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=73020 $Y=75670 $D=28
M1462 2212 2209 308 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.104e-13 pd=8e-07 ps=1.08e-06 nrd=0.166667 nrs=0.306667 sa=1.48017e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=73500 $Y=75550 $D=28
M1463 VSS 277 2212 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.48455e-13 as=6e-14 pd=2.03182e-06 ps=8e-07 nrd=0.690152 nrs=0.166667 sa=1.62933e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=73820 $Y=75550 $D=28
M1464 2214 761 2213 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=1.728e-13 pd=7.4e-07 ps=1.72e-06 nrd=0.185185 nrs=0.592593 sa=3.2e-07 sb=1.6437e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=179890 $Y=27120 $D=28
M1465 VSS 741 2214 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21728e-13 as=5.4e-14 pd=1.23972e-06 ps=7.4e-07 nrd=0.417449 nrs=0.185185 sa=6.4e-07 sb=1.54389e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=180210 $Y=27120 $D=28
M1466 2215 756 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.35254e-13 pd=8e-07 ps=1.37746e-06 nrd=0.166667 nrs=0.375704 sa=8.48167e-07 sb=1.288e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=180700 $Y=26930 $D=28
M1467 780 2213 2215 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.104e-13 as=6e-14 pd=1.08e-06 ps=8e-07 nrd=0.306667 nrs=0.166667 sa=1.16817e-06 sb=9.68e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=181020 $Y=26930 $D=28
M1468 2216 2213 780 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=1.104e-13 pd=8e-07 ps=1.08e-06 nrd=0.166667 nrs=0.306667 sa=1.48017e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=181500 $Y=27050 $D=28
M1469 VSS 756 2216 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.48455e-13 as=6e-14 pd=2.03182e-06 ps=8e-07 nrd=0.690152 nrs=0.166667 sa=1.62933e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=181820 $Y=27050 $D=28
M1470 2218 853 2217 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.28e-14 as=1.536e-13 pd=7e-07 ps=1.6e-06 nrd=0.229167 nrs=0.666667 sa=3.2e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=141670 $Y=27230 $D=28
M1471 VSS 536 2218 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3824e-13 as=5.28e-14 pd=9.80571e-07 ps=7e-07 nrd=0.6 nrs=0.229167 sa=6.6e-07 sb=9.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=142010 $Y=27230 $D=28
M1472 555 2217 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.6496e-13 pd=2.48e-06 ps=1.87943e-06 nrd=0.347826 nrs=0.313043 sa=8.45217e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=142640 $Y=26790 $D=28
M1473 2220 602 2219 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.28e-14 as=1.536e-13 pd=7e-07 ps=1.6e-06 nrd=0.229167 nrs=0.666667 sa=3.2e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=152470 $Y=63230 $D=28
M1474 VSS 614 2220 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3824e-13 as=5.28e-14 pd=9.80571e-07 ps=7e-07 nrd=0.6 nrs=0.229167 sa=6.6e-07 sb=9.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=152810 $Y=63230 $D=28
M1475 608 2219 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.6496e-13 pd=2.48e-06 ps=1.87943e-06 nrd=0.347826 nrs=0.313043 sa=8.45217e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=153440 $Y=62790 $D=28
M1476 2222 720 2221 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.28e-14 as=1.536e-13 pd=7e-07 ps=1.6e-06 nrd=0.229167 nrs=0.666667 sa=3.2e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=177270 $Y=39490 $D=28
M1477 VSS 735 2222 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3824e-13 as=5.28e-14 pd=9.80571e-07 ps=7e-07 nrd=0.6 nrs=0.229167 sa=6.6e-07 sb=9.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=177610 $Y=39490 $D=28
M1478 778 2221 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.6496e-13 pd=2.48e-06 ps=1.87943e-06 nrd=0.347826 nrs=0.313043 sa=8.45217e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=178240 $Y=39490 $D=28
M1479 2224 732 2223 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.28e-14 as=1.536e-13 pd=7e-07 ps=1.6e-06 nrd=0.229167 nrs=0.666667 sa=3.2e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=177670 $Y=56030 $D=28
M1480 VSS 734 2224 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3824e-13 as=5.28e-14 pd=9.80571e-07 ps=7e-07 nrd=0.6 nrs=0.229167 sa=6.6e-07 sb=9.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=178010 $Y=56030 $D=28
M1481 753 2223 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.6496e-13 pd=2.48e-06 ps=1.87943e-06 nrd=0.347826 nrs=0.313043 sa=8.45217e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=178640 $Y=55590 $D=28
M1482 2226 737 2225 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.28e-14 as=1.536e-13 pd=7e-07 ps=1.6e-06 nrd=0.229167 nrs=0.666667 sa=3.2e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=178470 $Y=25090 $D=28
M1483 VSS 761 2226 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3824e-13 as=5.28e-14 pd=9.80571e-07 ps=7e-07 nrd=0.6 nrs=0.229167 sa=6.6e-07 sb=9.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=178810 $Y=25090 $D=28
M1484 755 2225 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.6496e-13 pd=2.48e-06 ps=1.87943e-06 nrd=0.347826 nrs=0.313043 sa=8.45217e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=179440 $Y=25090 $D=28
M1485 VSS 666 2227 VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=1.28e-13 pd=7.6e-07 ps=1.44e-06 nrd=0.45 nrs=0.8 sa=3.2e-07 sb=1.12875e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.56e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=162840 $Y=54260 $D=28
M1486 2227 659 VSS VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.135e-14 as=7.2e-14 pd=8.7e-07 ps=7.6e-07 nrd=0.508437 nrs=0.45 sa=8e-07 sb=6.4875e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.56e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=163320 $Y=54260 $D=28
M1487 650 633 2227 VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28e-13 as=8.135e-14 pd=1.44e-06 ps=8.7e-07 nrd=0.8 nrs=0.508437 sa=1.005e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=163800 $Y=54150 $D=28
M1488 VSS 863 2229 VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=1.28e-13 pd=7.6e-07 ps=1.44e-06 nrd=0.45 nrs=0.8 sa=3.2e-07 sb=1.12875e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.56e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=174440 $Y=55740 $D=28
M1489 2229 725 VSS VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.135e-14 as=7.2e-14 pd=8.7e-07 ps=7.6e-07 nrd=0.508437 nrs=0.45 sa=8e-07 sb=6.4875e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.56e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=174920 $Y=55740 $D=28
M1490 718 714 2229 VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28e-13 as=8.135e-14 pd=1.44e-06 ps=8.7e-07 nrd=0.8 nrs=0.508437 sa=1.005e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=175400 $Y=55850 $D=28
M1491 VSS 713 2231 VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=1.28e-13 pd=7.6e-07 ps=1.44e-06 nrd=0.45 nrs=0.8 sa=3.2e-07 sb=1.12875e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.56e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=178040 $Y=54260 $D=28
M1492 2231 659 VSS VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.135e-14 as=7.2e-14 pd=8.7e-07 ps=7.6e-07 nrd=0.508437 nrs=0.45 sa=8e-07 sb=6.4875e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.56e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=178520 $Y=54260 $D=28
M1493 739 721 2231 VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28e-13 as=8.135e-14 pd=1.44e-06 ps=8.7e-07 nrd=0.8 nrs=0.508437 sa=1.005e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=179000 $Y=54150 $D=28
M1494 VSS clk 2233 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=9290 $Y=63260 $D=28
M1495 2235 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=9730 $Y=63320 $D=28
M1496 VSS 2233 2238 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=10950 $Y=63190 $D=28
M1497 2234 18 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=11470 $Y=63350 $D=28
M1498 2243 2235 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=12450 $Y=63110 $D=28
M1499 2236 2234 2243 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=12770 $Y=63110 $D=28
M1500 2245 2238 2236 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=13300 $Y=63570 $D=28
M1501 VSS 2237 2245 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=13620 $Y=63570 $D=28
M1502 2246 32 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=14040 $Y=62790 $D=28
M1503 2237 2236 2246 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=14360 $Y=62790 $D=28
M1504 2240 2238 2237 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=14840 $Y=63110 $D=28
M1505 2247 2235 2240 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=15420 $Y=63230 $D=28
M1506 2248 32 2247 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=15740 $Y=63230 $D=28
M1507 VSS 2239 2248 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=16060 $Y=63230 $D=28
M1508 VSS 2240 2239 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=17820 $Y=63510 $D=28
M1509 260 2240 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=18220 $Y=62790 $D=28
M1510 VSS clk 2250 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=96490 $Y=32400 $D=28
M1511 2252 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=96930 $Y=32400 $D=28
M1512 VSS 2250 2255 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=98150 $Y=32370 $D=28
M1513 2251 386 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=98670 $Y=32370 $D=28
M1514 2260 2252 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=99650 $Y=32150 $D=28
M1515 2253 2251 2260 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=99970 $Y=32150 $D=28
M1516 2262 2255 2253 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=100500 $Y=32230 $D=28
M1517 VSS 2254 2262 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=100820 $Y=32230 $D=28
M1518 2263 374 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=101240 $Y=32230 $D=28
M1519 2254 2253 2263 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=101560 $Y=32230 $D=28
M1520 2257 2255 2254 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=102040 $Y=32230 $D=28
M1521 2264 2252 2257 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=102620 $Y=32570 $D=28
M1522 2265 374 2264 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=102940 $Y=32570 $D=28
M1523 VSS 2256 2265 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=103260 $Y=32570 $D=28
M1524 VSS 2257 2256 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=105020 $Y=32290 $D=28
M1525 363 2257 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=105420 $Y=32290 $D=28
M1526 VSS clk 2267 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=109290 $Y=20060 $D=28
M1527 2269 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=109730 $Y=20120 $D=28
M1528 VSS 2267 2272 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=110950 $Y=19990 $D=28
M1529 2268 834 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=111470 $Y=20150 $D=28
M1530 2277 2269 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=112450 $Y=19910 $D=28
M1531 2270 2268 2277 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=112770 $Y=19910 $D=28
M1532 2279 2272 2270 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=113300 $Y=20370 $D=28
M1533 VSS 2271 2279 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=113620 $Y=20370 $D=28
M1534 2280 425 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=114040 $Y=19590 $D=28
M1535 2271 2270 2280 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=114360 $Y=19590 $D=28
M1536 2274 2272 2271 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=114840 $Y=19910 $D=28
M1537 2281 2269 2274 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=115420 $Y=20030 $D=28
M1538 2282 425 2281 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=115740 $Y=20030 $D=28
M1539 VSS 2273 2282 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=116060 $Y=20030 $D=28
M1540 VSS 2274 2273 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=117820 $Y=20310 $D=28
M1541 474 2274 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=118220 $Y=19590 $D=28
M1542 VSS clk 2284 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=119290 $Y=46800 $D=28
M1543 2286 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=119730 $Y=46800 $D=28
M1544 VSS 2284 2289 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=120950 $Y=46770 $D=28
M1545 2285 475 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=121470 $Y=46770 $D=28
M1546 2294 2286 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=122450 $Y=46550 $D=28
M1547 2287 2285 2294 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=122770 $Y=46550 $D=28
M1548 2296 2289 2287 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=123300 $Y=46630 $D=28
M1549 VSS 2288 2296 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=123620 $Y=46630 $D=28
M1550 2297 543 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=124040 $Y=46630 $D=28
M1551 2288 2287 2297 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=124360 $Y=46630 $D=28
M1552 2291 2289 2288 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=124840 $Y=46630 $D=28
M1553 2298 2286 2291 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=125420 $Y=46970 $D=28
M1554 2299 543 2298 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=125740 $Y=46970 $D=28
M1555 VSS 2290 2299 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=126060 $Y=46970 $D=28
M1556 VSS 2291 2290 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=127820 $Y=46690 $D=28
M1557 444 2291 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=128220 $Y=46690 $D=28
M1558 VSS clk 2301 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=134890 $Y=25200 $D=28
M1559 2303 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=135330 $Y=25200 $D=28
M1560 VSS 2301 2306 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=136550 $Y=25170 $D=28
M1561 2302 852 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=137070 $Y=25170 $D=28
M1562 2311 2303 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=138050 $Y=24950 $D=28
M1563 2304 2302 2311 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=138370 $Y=24950 $D=28
M1564 2313 2306 2304 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=138900 $Y=25030 $D=28
M1565 VSS 2305 2313 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=139220 $Y=25030 $D=28
M1566 2314 479 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=139640 $Y=25030 $D=28
M1567 2305 2304 2314 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=139960 $Y=25030 $D=28
M1568 2308 2306 2305 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=140440 $Y=25030 $D=28
M1569 2315 2303 2308 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=141020 $Y=25370 $D=28
M1570 2316 479 2315 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=141340 $Y=25370 $D=28
M1571 VSS 2307 2316 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=141660 $Y=25370 $D=28
M1572 VSS 2308 2307 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=143420 $Y=25090 $D=28
M1573 505 2308 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=143820 $Y=25090 $D=28
M1574 VSS clk 2318 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=146090 $Y=70460 $D=28
M1575 2320 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=146530 $Y=70520 $D=28
M1576 VSS 2318 2323 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=147750 $Y=70390 $D=28
M1577 2319 552 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=148270 $Y=70550 $D=28
M1578 2328 2320 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=149250 $Y=70310 $D=28
M1579 2321 2319 2328 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=149570 $Y=70310 $D=28
M1580 2330 2323 2321 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=150100 $Y=70770 $D=28
M1581 VSS 2322 2330 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=150420 $Y=70770 $D=28
M1582 2331 610 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=150840 $Y=69990 $D=28
M1583 2322 2321 2331 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=151160 $Y=69990 $D=28
M1584 2325 2323 2322 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=151640 $Y=70310 $D=28
M1585 2332 2320 2325 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=152220 $Y=70430 $D=28
M1586 2333 610 2332 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=152540 $Y=70430 $D=28
M1587 VSS 2324 2333 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=152860 $Y=70430 $D=28
M1588 VSS 2325 2324 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=154620 $Y=70710 $D=28
M1589 617 2325 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=155020 $Y=69990 $D=28
M1590 VSS clk 2335 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=149290 $Y=34460 $D=28
M1591 2337 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=149730 $Y=34520 $D=28
M1592 VSS 2335 2340 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=150950 $Y=34390 $D=28
M1593 2336 596 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=151470 $Y=34550 $D=28
M1594 2345 2337 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=152450 $Y=34310 $D=28
M1595 2338 2336 2345 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=152770 $Y=34310 $D=28
M1596 2347 2340 2338 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=153300 $Y=34770 $D=28
M1597 VSS 2339 2347 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=153620 $Y=34770 $D=28
M1598 2348 564 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=154040 $Y=33990 $D=28
M1599 2339 2338 2348 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=154360 $Y=33990 $D=28
M1600 2342 2340 2339 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=154840 $Y=34310 $D=28
M1601 2349 2337 2342 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=155420 $Y=34430 $D=28
M1602 2350 564 2349 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=155740 $Y=34430 $D=28
M1603 VSS 2341 2350 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=156060 $Y=34430 $D=28
M1604 VSS 2342 2341 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=157820 $Y=34710 $D=28
M1605 632 2342 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=158220 $Y=33990 $D=28
M1606 VSS clk 2352 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=150490 $Y=46800 $D=28
M1607 2354 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=150930 $Y=46800 $D=28
M1608 VSS 2352 2357 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=152150 $Y=46770 $D=28
M1609 2353 606 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=152670 $Y=46770 $D=28
M1610 2362 2354 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=153650 $Y=46550 $D=28
M1611 2355 2353 2362 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=153970 $Y=46550 $D=28
M1612 2364 2357 2355 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=154500 $Y=46630 $D=28
M1613 VSS 2356 2364 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=154820 $Y=46630 $D=28
M1614 2365 697 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=155240 $Y=46630 $D=28
M1615 2356 2355 2365 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=155560 $Y=46630 $D=28
M1616 2359 2357 2356 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=156040 $Y=46630 $D=28
M1617 2366 2354 2359 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=156620 $Y=46970 $D=28
M1618 2367 697 2366 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=156940 $Y=46970 $D=28
M1619 VSS 2358 2367 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=157260 $Y=46970 $D=28
M1620 VSS 2359 2358 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=159020 $Y=46690 $D=28
M1621 646 2359 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=159420 $Y=46690 $D=28
M1622 VSS clk 2369 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=156490 $Y=63260 $D=28
M1623 2371 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=156930 $Y=63320 $D=28
M1624 VSS 2369 2374 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=158150 $Y=63190 $D=28
M1625 2370 858 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=158670 $Y=63350 $D=28
M1626 2379 2371 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=159650 $Y=63110 $D=28
M1627 2372 2370 2379 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=159970 $Y=63110 $D=28
M1628 2381 2374 2372 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=160500 $Y=63570 $D=28
M1629 VSS 2373 2381 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=160820 $Y=63570 $D=28
M1630 2382 610 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=161240 $Y=62790 $D=28
M1631 2373 2372 2382 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=161560 $Y=62790 $D=28
M1632 2376 2374 2373 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=162040 $Y=63110 $D=28
M1633 2383 2371 2376 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=162620 $Y=63230 $D=28
M1634 2384 610 2383 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=162940 $Y=63230 $D=28
M1635 VSS 2375 2384 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=163260 $Y=63230 $D=28
M1636 VSS 2376 2375 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=165020 $Y=63510 $D=28
M1637 652 2376 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=165420 $Y=62790 $D=28
M1638 VSS clk 2386 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=159290 $Y=34460 $D=28
M1639 2388 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=159730 $Y=34520 $D=28
M1640 VSS 2386 2391 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=160950 $Y=34390 $D=28
M1641 2387 694 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=161470 $Y=34550 $D=28
M1642 2396 2388 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=162450 $Y=34310 $D=28
M1643 2389 2387 2396 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=162770 $Y=34310 $D=28
M1644 2398 2391 2389 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=163300 $Y=34770 $D=28
M1645 VSS 2390 2398 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=163620 $Y=34770 $D=28
M1646 2399 760 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=164040 $Y=33990 $D=28
M1647 2390 2389 2399 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=164360 $Y=33990 $D=28
M1648 2393 2391 2390 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=164840 $Y=34310 $D=28
M1649 2400 2388 2393 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=165420 $Y=34430 $D=28
M1650 2401 760 2400 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=165740 $Y=34430 $D=28
M1651 VSS 2392 2401 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=166060 $Y=34430 $D=28
M1652 VSS 2393 2392 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=167820 $Y=34710 $D=28
M1653 683 2393 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=168220 $Y=33990 $D=28
M1654 VSS clk 2403 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=164090 $Y=70460 $D=28
M1655 2405 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=164530 $Y=70520 $D=28
M1656 VSS 2403 2408 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=165750 $Y=70390 $D=28
M1657 2404 859 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=166270 $Y=70550 $D=28
M1658 2413 2405 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=167250 $Y=70310 $D=28
M1659 2406 2404 2413 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=167570 $Y=70310 $D=28
M1660 2415 2408 2406 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=168100 $Y=70770 $D=28
M1661 VSS 2407 2415 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=168420 $Y=70770 $D=28
M1662 2416 610 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=168840 $Y=69990 $D=28
M1663 2407 2406 2416 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=169160 $Y=69990 $D=28
M1664 2410 2408 2407 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=169640 $Y=70310 $D=28
M1665 2417 2405 2410 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=170220 $Y=70430 $D=28
M1666 2418 610 2417 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=170540 $Y=70430 $D=28
M1667 VSS 2409 2418 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=170860 $Y=70430 $D=28
M1668 VSS 2410 2409 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=172620 $Y=70710 $D=28
M1669 576 2410 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=173020 $Y=69990 $D=28
M1670 VSS clk 2420 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=169690 $Y=27260 $D=28
M1671 2422 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=170130 $Y=27320 $D=28
M1672 VSS 2420 2425 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=171350 $Y=27190 $D=28
M1673 2421 704 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=171870 $Y=27350 $D=28
M1674 2430 2422 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=172850 $Y=27110 $D=28
M1675 2423 2421 2430 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=173170 $Y=27110 $D=28
M1676 2432 2425 2423 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=173700 $Y=27570 $D=28
M1677 VSS 2424 2432 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=174020 $Y=27570 $D=28
M1678 2433 706 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=174440 $Y=26790 $D=28
M1679 2424 2423 2433 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=174760 $Y=26790 $D=28
M1680 2427 2425 2424 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=175240 $Y=27110 $D=28
M1681 2434 2422 2427 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=175820 $Y=27230 $D=28
M1682 2435 706 2434 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=176140 $Y=27230 $D=28
M1683 VSS 2426 2435 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=176460 $Y=27230 $D=28
M1684 VSS 2427 2426 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=178220 $Y=27510 $D=28
M1685 716 2427 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=178620 $Y=26790 $D=28
M1686 VSS clk 2437 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=175690 $Y=12860 $D=28
M1687 2439 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=176130 $Y=12920 $D=28
M1688 VSS 2437 2442 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=177350 $Y=12790 $D=28
M1689 2438 754 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=177870 $Y=12950 $D=28
M1690 2447 2439 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=178850 $Y=12710 $D=28
M1691 2440 2438 2447 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=179170 $Y=12710 $D=28
M1692 2449 2442 2440 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=179700 $Y=13170 $D=28
M1693 VSS 2441 2449 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=180020 $Y=13170 $D=28
M1694 2450 706 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=180440 $Y=12390 $D=28
M1695 2441 2440 2450 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=180760 $Y=12390 $D=28
M1696 2444 2442 2441 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=181240 $Y=12710 $D=28
M1697 2451 2439 2444 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=181820 $Y=12830 $D=28
M1698 2452 706 2451 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=182140 $Y=12830 $D=28
M1699 VSS 2443 2452 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=182460 $Y=12830 $D=28
M1700 VSS 2444 2443 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=184220 $Y=13110 $D=28
M1701 733 2444 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=184620 $Y=12390 $D=28
M1702 VSS clk 2454 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=175690 $Y=68400 $D=28
M1703 2456 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=176130 $Y=68400 $D=28
M1704 VSS 2454 2459 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=177350 $Y=68370 $D=28
M1705 2455 762 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=177870 $Y=68370 $D=28
M1706 2464 2456 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=178850 $Y=68150 $D=28
M1707 2457 2455 2464 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=179170 $Y=68150 $D=28
M1708 2466 2459 2457 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=179700 $Y=68230 $D=28
M1709 VSS 2458 2466 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=180020 $Y=68230 $D=28
M1710 2467 760 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=180440 $Y=68230 $D=28
M1711 2458 2457 2467 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=180760 $Y=68230 $D=28
M1712 2461 2459 2458 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=181240 $Y=68230 $D=28
M1713 2468 2456 2461 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=181820 $Y=68570 $D=28
M1714 2469 760 2468 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=182140 $Y=68570 $D=28
M1715 VSS 2460 2469 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=182460 $Y=68570 $D=28
M1716 VSS 2461 2460 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=184220 $Y=68290 $D=28
M1717 746 2461 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=184620 $Y=68290 $D=28
M1718 VSS clk 2471 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=176090 $Y=34460 $D=28
M1719 2473 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=176530 $Y=34520 $D=28
M1720 VSS 2471 2476 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=177750 $Y=34390 $D=28
M1721 2472 782 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=178270 $Y=34550 $D=28
M1722 2481 2473 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=179250 $Y=34310 $D=28
M1723 2474 2472 2481 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=179570 $Y=34310 $D=28
M1724 2483 2476 2474 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=180100 $Y=34770 $D=28
M1725 VSS 2475 2483 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=180420 $Y=34770 $D=28
M1726 2484 706 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=180840 $Y=33990 $D=28
M1727 2475 2474 2484 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=181160 $Y=33990 $D=28
M1728 2478 2476 2475 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=181640 $Y=34310 $D=28
M1729 2485 2473 2478 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=182220 $Y=34430 $D=28
M1730 2486 706 2485 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=182540 $Y=34430 $D=28
M1731 VSS 2477 2486 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=182860 $Y=34430 $D=28
M1732 VSS 2478 2477 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=184620 $Y=34710 $D=28
M1733 717 2478 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=185020 $Y=33990 $D=28
M1734 VSS clk 2488 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.54581e-14 as=1.088e-13 pd=8.99355e-07 ps=1.32e-06 nrd=0.652751 nrs=0.941176 sa=3.2e-07 sb=7.17647e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.8e-14 panw8=0 panw9=0 panw10=0 $X=177690 $Y=48860 $D=28
M1735 2490 clk VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.064e-13 as=6.21419e-14 pd=1.32e-06 ps=7.40645e-07 nrd=1.35714 nrs=0.792627 sa=7.6e-07 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=4.8e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=178130 $Y=48920 $D=28
M1736 VSS 2488 2493 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.39523e-13 as=1.408e-13 pd=1.27032e-06 ps=1.52e-06 nrd=0.720674 nrs=0.727273 sa=3.2e-07 sb=6.50909e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=179350 $Y=48790 $D=28
M1737 2489 864 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.87871e-14 pd=1.2e-06 ps=8.08387e-07 nrd=1.14286 nrs=1.13249 sa=8.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=179870 $Y=48950 $D=28
M1738 2498 2490 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4e-14 as=2.34652e-13 pd=9.4e-07 ps=2.13645e-06 nrd=0.135135 nrs=0.428509 sa=3.6e-07 sb=1.00649e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=180850 $Y=48710 $D=28
M1739 2491 2489 2498 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.99957e-13 as=7.4e-14 pd=1.81064e-06 ps=9.4e-07 nrd=0.365152 nrs=0.135135 sa=6.8e-07 sb=7.72973e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=181170 $Y=48710 $D=28
M1740 2500 2493 2491 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.40426e-14 pd=4e-07 ps=4.89362e-07 nrd=0.5 nrs=1.35106 sa=1.21e-06 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=181700 $Y=49170 $D=28
M1741 VSS 2492 2500 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.25753e-14 as=2e-14 pd=4.68493e-07 ps=4e-07 nrd=1.06438 nrs=0.5 sa=1.53e-06 sb=1.54e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=182020 $Y=49170 $D=28
M1742 2501 760 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.08619e-13 pd=1.18e-06 ps=2.29562e-06 nrd=0.102041 nrs=0.217221 sa=5.76735e-07 sb=1.1098e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=182440 $Y=48390 $D=28
M1743 2492 2491 2501 VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80224e-13 as=9.8e-14 pd=1.60146e-06 ps=1.18e-06 nrd=0.187656 nrs=0.102041 sa=8.41633e-07 sb=8.55102e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=182760 $Y=48390 $D=28
M1744 2495 2493 2492 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.88177e-13 as=1.21376e-13 pd=1.71907e-06 ps=1.07854e-06 nrd=0.431994 nrs=0.27864 sa=1.30303e-06 sb=7.1697e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=183240 $Y=48710 $D=28
M1745 2502 2490 2495 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=5.70233e-14 pd=4e-07 ps=5.2093e-07 nrd=0.5 nrs=1.42558 sa=1.58e-06 sb=1.02e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=183820 $Y=48830 $D=28
M1746 2503 760 2502 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.9e-06 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=184140 $Y=48830 $D=28
M1747 VSS 2494 2503 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09833e-13 as=2e-14 pd=1.04167e-06 ps=4e-07 nrd=2.74583 nrs=0.5 sa=2e-06 sb=3.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=9.6e-15 panw8=1.44e-14 panw9=0 panw10=0 $X=184460 $Y=48830 $D=28
M1748 VSS 2495 2494 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.17143e-14 as=1.056e-13 pd=4.71429e-07 ps=1.36e-06 nrd=1.04286 nrs=2.64 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=186220 $Y=49110 $D=28
M1749 726 2495 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.22e-13 as=1.91886e-13 pd=2.54e-06 ps=2.16857e-06 nrd=0.380435 nrs=0.226708 sa=3.58261e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=186620 $Y=48390 $D=28
M1750 2507 256 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=70070 $Y=13050 $D=28
M1751 2506 264 2507 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=70390 $Y=13050 $D=28
M1752 2508 310 2506 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=70960 $Y=13050 $D=28
M1753 VSS result[1] 2508 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=71280 $Y=13050 $D=28
M1754 251 2506 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=71830 $Y=13070 $D=28
M1755 2511 256 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=76470 $Y=13050 $D=28
M1756 2510 143 2511 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=76790 $Y=13050 $D=28
M1757 2512 310 2510 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=77360 $Y=13050 $D=28
M1758 VSS result[2] 2512 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=77680 $Y=13050 $D=28
M1759 828 2510 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=78230 $Y=13070 $D=28
M1760 2515 256 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=79270 $Y=13050 $D=28
M1761 2514 298 2515 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=79590 $Y=13050 $D=28
M1762 2516 310 2514 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=80160 $Y=13050 $D=28
M1763 VSS result[0] 2516 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=80480 $Y=13050 $D=28
M1764 269 2514 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=81030 $Y=13070 $D=28
M1765 2519 300 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=80070 $Y=32290 $D=28
M1766 2518 159 2519 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=80390 $Y=32290 $D=28
M1767 2520 306 2518 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=80960 $Y=32290 $D=28
M1768 VSS result[5] 2520 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=81280 $Y=32290 $D=28
M1769 305 2518 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=81830 $Y=32290 $D=28
M1770 2523 300 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=82870 $Y=32290 $D=28
M1771 2522 109 2523 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=83190 $Y=32290 $D=28
M1772 2524 306 2522 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=83760 $Y=32290 $D=28
M1773 VSS result[6] 2524 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=84080 $Y=32290 $D=28
M1774 321 2522 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=84630 $Y=32290 $D=28
M1775 2527 318 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=85670 $Y=20250 $D=28
M1776 2526 62 2527 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=85990 $Y=20250 $D=28
M1777 2528 345 2526 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=86560 $Y=20250 $D=28
M1778 VSS result[4] 2528 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=86880 $Y=20250 $D=28
M1779 322 2526 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=87430 $Y=20270 $D=28
M1780 2531 389 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=88470 $Y=13050 $D=28
M1781 2530 100 2531 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=88790 $Y=13050 $D=28
M1782 2532 326 2530 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=89360 $Y=13050 $D=28
M1783 VSS result[3] 2532 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=89680 $Y=13050 $D=28
M1784 333 2530 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=90230 $Y=13070 $D=28
M1785 2535 318 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=88870 $Y=20250 $D=28
M1786 2534 260 2535 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=89190 $Y=20250 $D=28
M1787 2536 345 2534 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=89760 $Y=20250 $D=28
M1788 VSS result[7] 2536 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=90080 $Y=20250 $D=28
M1789 332 2534 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=90630 $Y=20270 $D=28
M1790 2539 377 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96070 $Y=20250 $D=28
M1791 2538 239 2539 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96390 $Y=20250 $D=28
M1792 2540 368 2538 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96960 $Y=20250 $D=28
M1793 VSS result[8] 2540 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=97280 $Y=20250 $D=28
M1794 832 2538 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=97830 $Y=20270 $D=28
M1795 2543 389 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=97270 $Y=13050 $D=28
M1796 2542 359 2543 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=97590 $Y=13050 $D=28
M1797 2544 326 2542 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=98160 $Y=13050 $D=28
M1798 VSS result[10] 2544 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=98480 $Y=13050 $D=28
M1799 364 2542 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=99030 $Y=13070 $D=28
M1800 2547 399 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=100070 $Y=20250 $D=28
M1801 2546 363 2547 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=100390 $Y=20250 $D=28
M1802 2548 368 2546 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=100960 $Y=20250 $D=28
M1803 VSS result[9] 2548 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=101280 $Y=20250 $D=28
M1804 373 2546 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=101830 $Y=20270 $D=28
M1805 2551 389 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=102470 $Y=13050 $D=28
M1806 2550 418 2551 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=102790 $Y=13050 $D=28
M1807 2552 326 2550 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=103360 $Y=13050 $D=28
M1808 VSS result[11] 2552 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=103680 $Y=13050 $D=28
M1809 385 2550 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=104230 $Y=13070 $D=28
M1810 2555 408 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=106870 $Y=17890 $D=28
M1811 2554 452 2555 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=107190 $Y=17890 $D=28
M1812 2556 396 2554 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=107760 $Y=17890 $D=28
M1813 VSS result[12] 2556 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=108080 $Y=17890 $D=28
M1814 388 2554 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=108630 $Y=17890 $D=28
M1815 2559 408 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=118870 $Y=17890 $D=28
M1816 2558 444 2559 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=119190 $Y=17890 $D=28
M1817 2560 396 2558 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=119760 $Y=17890 $D=28
M1818 VSS result[14] 2560 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=120080 $Y=17890 $D=28
M1819 453 2558 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=120630 $Y=17890 $D=28
M1820 2563 408 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=118870 $Y=25090 $D=28
M1821 2562 839 2563 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=119190 $Y=25090 $D=28
M1822 2564 396 2562 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=119760 $Y=25090 $D=28
M1823 VSS result[13] 2564 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=120080 $Y=25090 $D=28
M1824 454 2562 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=120630 $Y=25090 $D=28
M1825 2567 491 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=123670 $Y=13050 $D=28
M1826 2566 456 2567 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=123990 $Y=13050 $D=28
M1827 2568 526 2566 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=124560 $Y=13050 $D=28
M1828 VSS result[15] 2568 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=124880 $Y=13050 $D=28
M1829 424 2566 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=125430 $Y=13070 $D=28
M1830 2571 491 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=126470 $Y=13050 $D=28
M1831 2570 474 2571 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=126790 $Y=13050 $D=28
M1832 2572 526 2570 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=127360 $Y=13050 $D=28
M1833 VSS result[16] 2572 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=127680 $Y=13050 $D=28
M1834 449 2570 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=128230 $Y=13070 $D=28
M1835 2575 500 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=131270 $Y=13050 $D=28
M1836 2574 505 2575 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=131590 $Y=13050 $D=28
M1837 2576 526 2574 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=132160 $Y=13050 $D=28
M1838 VSS result[17] 2576 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=132480 $Y=13050 $D=28
M1839 513 2574 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=133030 $Y=13070 $D=28
M1840 2579 500 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=136870 $Y=13050 $D=28
M1841 2578 568 2579 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=137190 $Y=13050 $D=28
M1842 2580 570 2578 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=137760 $Y=13050 $D=28
M1843 VSS result[18] 2580 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=138080 $Y=13050 $D=28
M1844 541 2578 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=138630 $Y=13070 $D=28
M1845 2583 611 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=145270 $Y=17890 $D=28
M1846 2582 632 2583 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=145590 $Y=17890 $D=28
M1847 2584 570 2582 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=146160 $Y=17890 $D=28
M1848 VSS result[19] 2584 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=146480 $Y=17890 $D=28
M1849 579 2582 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=147030 $Y=17890 $D=28
M1850 2587 593 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=150470 $Y=17890 $D=28
M1851 2586 597 2587 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=150790 $Y=17890 $D=28
M1852 2588 620 2586 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=151360 $Y=17890 $D=28
M1853 VSS result[21] 2588 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=151680 $Y=17890 $D=28
M1854 604 2586 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=152230 $Y=17890 $D=28
M1855 2591 593 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=154870 $Y=17890 $D=28
M1856 2590 646 2591 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=155190 $Y=17890 $D=28
M1857 2592 570 2590 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=155760 $Y=17890 $D=28
M1858 VSS result[20] 2592 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=156080 $Y=17890 $D=28
M1859 623 2590 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=156630 $Y=17890 $D=28
M1860 2595 688 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=156470 $Y=32290 $D=28
M1861 2594 652 2595 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=156790 $Y=32290 $D=28
M1862 2596 651 2594 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=157360 $Y=32290 $D=28
M1863 VSS result[25] 2596 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=157680 $Y=32290 $D=28
M1864 612 2594 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=158230 $Y=32290 $D=28
M1865 2599 593 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=157670 $Y=17890 $D=28
M1866 2598 609 2599 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=157990 $Y=17890 $D=28
M1867 2600 645 2598 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=158560 $Y=17890 $D=28
M1868 VSS result[22] 2600 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=158880 $Y=17890 $D=28
M1869 621 2598 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=159430 $Y=17890 $D=28
M1870 2603 682 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=157670 $Y=25090 $D=28
M1871 2602 576 2603 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=157990 $Y=25090 $D=28
M1872 2604 620 2602 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=158560 $Y=25090 $D=28
M1873 VSS result[24] 2604 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=158880 $Y=25090 $D=28
M1874 563 2602 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=159430 $Y=25090 $D=28
M1875 2607 682 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=160470 $Y=25090 $D=28
M1876 2606 617 2607 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=160790 $Y=25090 $D=28
M1877 2608 620 2606 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=161360 $Y=25090 $D=28
M1878 VSS result[23] 2608 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=161680 $Y=25090 $D=28
M1879 654 2606 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=162230 $Y=25090 $D=28
M1880 2611 689 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=161670 $Y=32290 $D=28
M1881 2610 746 2611 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=161990 $Y=32290 $D=28
M1882 2612 651 2610 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=162560 $Y=32290 $D=28
M1883 VSS result[26] 2612 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=162880 $Y=32290 $D=28
M1884 656 2610 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=163430 $Y=32290 $D=28
M1885 2615 688 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=164870 $Y=17890 $D=28
M1886 2614 683 2615 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=165190 $Y=17890 $D=28
M1887 2616 701 2614 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=165760 $Y=17890 $D=28
M1888 VSS result[28] 2616 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=166080 $Y=17890 $D=28
M1889 643 2614 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=166630 $Y=17890 $D=28
M1890 2619 682 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=166470 $Y=25090 $D=28
M1891 2618 726 2619 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=166790 $Y=25090 $D=28
M1892 2620 651 2618 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=167360 $Y=25090 $D=28
M1893 VSS result[27] 2620 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=167680 $Y=25090 $D=28
M1894 678 2618 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=168230 $Y=25090 $D=28
M1895 2623 688 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=170070 $Y=13050 $D=28
M1896 2622 717 2623 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=170390 $Y=13050 $D=28
M1897 2624 701 2622 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=170960 $Y=13050 $D=28
M1898 VSS result[29] 2624 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=171280 $Y=13050 $D=28
M1899 699 2622 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=171830 $Y=13070 $D=28
M1900 2627 693 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=172870 $Y=13050 $D=28
M1901 2626 716 2627 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=173190 $Y=13050 $D=28
M1902 2628 701 2626 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=173760 $Y=13050 $D=28
M1903 VSS result[30] 2628 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=174080 $Y=13050 $D=28
M1904 708 2626 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=174630 $Y=13070 $D=28
M1905 2631 693 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=2.668e-13 pd=4.6e-07 ps=2.48e-06 nrd=0.384615 nrs=3.94675 sa=3.8e-07 sb=1.96538e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=177270 $Y=17890 $D=28
M1906 2630 733 2631 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13e-14 as=2.6e-14 pd=7.3e-07 ps=4.6e-07 nrd=0.906805 nrs=0.384615 sa=7e-07 sb=1.75615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=177590 $Y=17890 $D=28
M1907 2632 701 2630 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.6e-14 as=6.13e-14 pd=4.6e-07 ps=7.3e-07 nrd=0.384615 nrs=0.906805 sa=1.27e-06 sb=1.18615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=178160 $Y=17890 $D=28
M1908 VSS result[31] 2632 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20933e-13 as=2.6e-14 pd=1.09333e-06 ps=4.6e-07 nrd=1.78895 nrs=0.384615 sa=1.59e-06 sb=8.66154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=178480 $Y=17890 $D=28
M1909 740 2630 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.11631e-13 pd=1.28e-06 ps=1.00923e-06 nrd=1.69444 nrs=1.93803 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=179030 $Y=17890 $D=28
M1910 2640 2633 2634 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=25660 $Y=13090 $D=28
M1911 2642 78 2640 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=25980 $Y=13090 $D=28
M1912 VSS 68 2642 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=26300 $Y=13090 $D=28
M1913 VSS clk 2633 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=27280 $Y=12840 $D=28
M1914 2636 2633 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=27790 $Y=12940 $D=28
M1915 2644 2636 2634 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=28810 $Y=13010 $D=28
M1916 2645 2635 2644 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=29130 $Y=13010 $D=28
M1917 VSS 68 2645 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=29450 $Y=13010 $D=28
M1918 2635 2634 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=29910 $Y=12870 $D=28
M1919 2637 2636 2635 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=30470 $Y=12870 $D=28
M1920 2647 2633 2637 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=31030 $Y=13110 $D=28
M1921 VSS 2639 2647 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=31350 $Y=13110 $D=28
M1922 2648 68 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=31790 $Y=13090 $D=28
M1923 2639 2637 2648 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=32110 $Y=13090 $D=28
M1924 2638 2639 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=32430 $Y=12390 $D=28
M1925 VSS 2638 919 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=33330 $Y=13070 $D=28
M1926 weight_out[3] 2639 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=33830 $Y=13070 $D=28
M1927 2656 2649 2650 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=72060 $Y=17910 $D=28
M1928 2658 269 2656 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=72380 $Y=17910 $D=28
M1929 VSS 316 2658 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=72700 $Y=17910 $D=28
M1930 VSS clk 2649 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=73680 $Y=18060 $D=28
M1931 2652 2649 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=74190 $Y=18060 $D=28
M1932 2660 2652 2650 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=75210 $Y=17990 $D=28
M1933 2661 2651 2660 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=75530 $Y=17990 $D=28
M1934 VSS 316 2661 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=75850 $Y=17990 $D=28
M1935 2651 2650 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=76310 $Y=18130 $D=28
M1936 2653 2652 2651 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=76870 $Y=18130 $D=28
M1937 2663 2649 2653 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=77430 $Y=17890 $D=28
M1938 VSS 2655 2663 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=77750 $Y=17890 $D=28
M1939 2664 316 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=78190 $Y=17890 $D=28
M1940 2655 2653 2664 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=78510 $Y=17890 $D=28
M1941 2654 2655 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=78830 $Y=18610 $D=28
M1942 VSS 2654 920 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=79730 $Y=17890 $D=28
M1943 result[0] 2655 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=80230 $Y=17890 $D=28
M1944 2672 2665 2666 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=82060 $Y=17910 $D=28
M1945 2674 322 2672 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=82380 $Y=17910 $D=28
M1946 VSS 316 2674 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=82700 $Y=17910 $D=28
M1947 VSS clk 2665 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=83680 $Y=18060 $D=28
M1948 2668 2665 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=84190 $Y=18060 $D=28
M1949 2676 2668 2666 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=85210 $Y=17990 $D=28
M1950 2677 2667 2676 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=85530 $Y=17990 $D=28
M1951 VSS 316 2677 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=85850 $Y=17990 $D=28
M1952 2667 2666 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=86310 $Y=18130 $D=28
M1953 2669 2668 2667 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=86870 $Y=18130 $D=28
M1954 2679 2665 2669 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=87430 $Y=17890 $D=28
M1955 VSS 2671 2679 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=87750 $Y=17890 $D=28
M1956 2680 316 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=88190 $Y=17890 $D=28
M1957 2671 2669 2680 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=88510 $Y=17890 $D=28
M1958 2670 2671 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=88830 $Y=18610 $D=28
M1959 VSS 2670 921 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=89730 $Y=17890 $D=28
M1960 result[4] 2671 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=90230 $Y=17890 $D=28
M1961 2688 2681 2682 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=87260 $Y=32310 $D=28
M1962 2690 321 2688 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=87580 $Y=32310 $D=28
M1963 VSS 303 2690 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=87900 $Y=32310 $D=28
M1964 VSS clk 2681 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=88880 $Y=32460 $D=28
M1965 2684 2681 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=89390 $Y=32460 $D=28
M1966 2692 2684 2682 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=90410 $Y=32390 $D=28
M1967 2693 2683 2692 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=90730 $Y=32390 $D=28
M1968 VSS 303 2693 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=91050 $Y=32390 $D=28
M1969 2683 2682 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=91510 $Y=32530 $D=28
M1970 2685 2684 2683 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=92070 $Y=32530 $D=28
M1971 2695 2681 2685 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=92630 $Y=32290 $D=28
M1972 VSS 2687 2695 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=92950 $Y=32290 $D=28
M1973 2696 303 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=93390 $Y=32290 $D=28
M1974 2687 2685 2696 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=93710 $Y=32290 $D=28
M1975 2686 2687 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=94030 $Y=33010 $D=28
M1976 VSS 2686 922 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=94930 $Y=32290 $D=28
M1977 result[6] 2687 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=95430 $Y=32290 $D=28
M1978 2704 2697 2698 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=95660 $Y=34690 $D=28
M1979 2706 192 2704 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=95980 $Y=34690 $D=28
M1980 VSS 374 2706 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96300 $Y=34690 $D=28
M1981 VSS clk 2697 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=97280 $Y=34440 $D=28
M1982 2700 2697 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=97790 $Y=34540 $D=28
M1983 2708 2700 2698 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=98810 $Y=34610 $D=28
M1984 2709 2699 2708 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=99130 $Y=34610 $D=28
M1985 VSS 374 2709 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=99450 $Y=34610 $D=28
M1986 2699 2698 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=99910 $Y=34470 $D=28
M1987 2701 2700 2699 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=100470 $Y=34470 $D=28
M1988 2711 2697 2701 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=101030 $Y=34710 $D=28
M1989 VSS 2703 2711 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=101350 $Y=34710 $D=28
M1990 2712 374 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=101790 $Y=34690 $D=28
M1991 2703 2701 2712 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=102110 $Y=34690 $D=28
M1992 2702 2703 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=102430 $Y=33990 $D=28
M1993 VSS 2702 923 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=103330 $Y=34670 $D=28
M1994 data_out[3] 2703 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=103830 $Y=34670 $D=28
M1995 2720 2713 2714 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96060 $Y=17910 $D=28
M1996 2722 373 2720 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96380 $Y=17910 $D=28
M1997 VSS 371 2722 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96700 $Y=17910 $D=28
M1998 VSS clk 2713 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=97680 $Y=18060 $D=28
M1999 2716 2713 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=98190 $Y=18060 $D=28
M2000 2724 2716 2714 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=99210 $Y=17990 $D=28
M2001 2725 2715 2724 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=99530 $Y=17990 $D=28
M2002 VSS 371 2725 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=99850 $Y=17990 $D=28
M2003 2715 2714 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=100310 $Y=18130 $D=28
M2004 2717 2716 2715 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=100870 $Y=18130 $D=28
M2005 2727 2713 2717 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=101430 $Y=17890 $D=28
M2006 VSS 2719 2727 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=101750 $Y=17890 $D=28
M2007 2728 371 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=102190 $Y=17890 $D=28
M2008 2719 2717 2728 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=102510 $Y=17890 $D=28
M2009 2718 2719 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=102830 $Y=18610 $D=28
M2010 VSS 2718 924 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=103730 $Y=17890 $D=28
M2011 result[9] 2719 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=104230 $Y=17890 $D=28
M2012 2736 2729 2730 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=101660 $Y=27490 $D=28
M2013 2738 254 2736 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=101980 $Y=27490 $D=28
M2014 VSS 374 2738 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=102300 $Y=27490 $D=28
M2015 VSS clk 2729 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=103280 $Y=27240 $D=28
M2016 2732 2729 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=103790 $Y=27340 $D=28
M2017 2740 2732 2730 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=104810 $Y=27410 $D=28
M2018 2741 2731 2740 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=105130 $Y=27410 $D=28
M2019 VSS 374 2741 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=105450 $Y=27410 $D=28
M2020 2731 2730 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=105910 $Y=27270 $D=28
M2021 2733 2732 2731 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=106470 $Y=27270 $D=28
M2022 2743 2729 2733 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=107030 $Y=27510 $D=28
M2023 VSS 2735 2743 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=107350 $Y=27510 $D=28
M2024 2744 374 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=107790 $Y=27490 $D=28
M2025 2735 2733 2744 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=108110 $Y=27490 $D=28
M2026 2734 2735 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=108430 $Y=26790 $D=28
M2027 VSS 2734 925 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=109330 $Y=27470 $D=28
M2028 data_out[2] 2735 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=109830 $Y=27470 $D=28
M2029 2752 2745 2746 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=105660 $Y=10710 $D=28
M2030 2754 385 2752 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=105980 $Y=10710 $D=28
M2031 VSS 371 2754 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=106300 $Y=10710 $D=28
M2032 VSS clk 2745 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=107280 $Y=10860 $D=28
M2033 2748 2745 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=107790 $Y=10860 $D=28
M2034 2756 2748 2746 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=108810 $Y=10790 $D=28
M2035 2757 2747 2756 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=109130 $Y=10790 $D=28
M2036 VSS 371 2757 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=109450 $Y=10790 $D=28
M2037 2747 2746 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=109910 $Y=10930 $D=28
M2038 2749 2748 2747 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=110470 $Y=10930 $D=28
M2039 2759 2745 2749 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=111030 $Y=10690 $D=28
M2040 VSS 2751 2759 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=111350 $Y=10690 $D=28
M2041 2760 371 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=111790 $Y=10690 $D=28
M2042 2751 2749 2760 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=112110 $Y=10690 $D=28
M2043 2750 2751 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=112430 $Y=11410 $D=28
M2044 VSS 2750 926 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=113330 $Y=10690 $D=28
M2045 result[11] 2751 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=113830 $Y=10690 $D=28
M2046 2768 2761 2762 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=109660 $Y=17910 $D=28
M2047 2770 454 2768 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=109980 $Y=17910 $D=28
M2048 VSS 428 2770 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=110300 $Y=17910 $D=28
M2049 VSS clk 2761 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=111280 $Y=18060 $D=28
M2050 2764 2761 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=111790 $Y=18060 $D=28
M2051 2772 2764 2762 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=112810 $Y=17990 $D=28
M2052 2773 2763 2772 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=113130 $Y=17990 $D=28
M2053 VSS 428 2773 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=113450 $Y=17990 $D=28
M2054 2763 2762 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=113910 $Y=18130 $D=28
M2055 2765 2764 2763 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=114470 $Y=18130 $D=28
M2056 2775 2761 2765 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=115030 $Y=17890 $D=28
M2057 VSS 2767 2775 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=115350 $Y=17890 $D=28
M2058 2776 428 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=115790 $Y=17890 $D=28
M2059 2767 2765 2776 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=116110 $Y=17890 $D=28
M2060 2766 2767 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=116430 $Y=18610 $D=28
M2061 VSS 2766 927 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=117330 $Y=17890 $D=28
M2062 result[13] 2767 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=117830 $Y=17890 $D=28
M2063 2784 2777 2778 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=109660 $Y=25110 $D=28
M2064 2786 287 2784 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=109980 $Y=25110 $D=28
M2065 VSS 407 2786 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=110300 $Y=25110 $D=28
M2066 VSS clk 2777 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=111280 $Y=25260 $D=28
M2067 2780 2777 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=111790 $Y=25260 $D=28
M2068 2788 2780 2778 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=112810 $Y=25190 $D=28
M2069 2789 2779 2788 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=113130 $Y=25190 $D=28
M2070 VSS 407 2789 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=113450 $Y=25190 $D=28
M2071 2779 2778 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=113910 $Y=25330 $D=28
M2072 2781 2780 2779 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=114470 $Y=25330 $D=28
M2073 2791 2777 2781 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=115030 $Y=25090 $D=28
M2074 VSS 2783 2791 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=115350 $Y=25090 $D=28
M2075 2792 407 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=115790 $Y=25090 $D=28
M2076 2783 2781 2792 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=116110 $Y=25090 $D=28
M2077 2782 2783 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=116430 $Y=25810 $D=28
M2078 VSS 2782 928 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=117330 $Y=25090 $D=28
M2079 data_out[1] 2783 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=117830 $Y=25090 $D=28
M2080 2800 2793 2794 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=110060 $Y=49090 $D=28
M2081 2802 494 2800 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=110380 $Y=49090 $D=28
M2082 VSS 425 2802 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=110700 $Y=49090 $D=28
M2083 VSS clk 2793 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=111680 $Y=48840 $D=28
M2084 2796 2793 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=112190 $Y=48940 $D=28
M2085 2804 2796 2794 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=113210 $Y=49010 $D=28
M2086 2805 2795 2804 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=113530 $Y=49010 $D=28
M2087 VSS 425 2805 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=113850 $Y=49010 $D=28
M2088 2795 2794 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=114310 $Y=48870 $D=28
M2089 2797 2796 2795 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=114870 $Y=48870 $D=28
M2090 2807 2793 2797 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=115430 $Y=49110 $D=28
M2091 VSS 2799 2807 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=115750 $Y=49110 $D=28
M2092 2808 425 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=116190 $Y=49090 $D=28
M2093 2799 2797 2808 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=116510 $Y=49090 $D=28
M2094 2798 2799 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=116830 $Y=48390 $D=28
M2095 VSS 2798 436 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=117730 $Y=49070 $D=28
M2096 839 2799 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=118230 $Y=49070 $D=28
M2097 2816 2809 2810 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=119260 $Y=20290 $D=28
M2098 2818 453 2816 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=119580 $Y=20290 $D=28
M2099 VSS 428 2818 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=119900 $Y=20290 $D=28
M2100 VSS clk 2809 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=120880 $Y=20040 $D=28
M2101 2812 2809 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=121390 $Y=20140 $D=28
M2102 2820 2812 2810 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=122410 $Y=20210 $D=28
M2103 2821 2811 2820 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=122730 $Y=20210 $D=28
M2104 VSS 428 2821 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=123050 $Y=20210 $D=28
M2105 2811 2810 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=123510 $Y=20070 $D=28
M2106 2813 2812 2811 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=124070 $Y=20070 $D=28
M2107 2823 2809 2813 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=124630 $Y=20310 $D=28
M2108 VSS 2815 2823 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=124950 $Y=20310 $D=28
M2109 2824 428 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=125390 $Y=20290 $D=28
M2110 2815 2813 2824 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=125710 $Y=20290 $D=28
M2111 2814 2815 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=126030 $Y=19590 $D=28
M2112 VSS 2814 929 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=126930 $Y=20270 $D=28
M2113 result[14] 2815 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=127430 $Y=20270 $D=28
M2114 2832 2825 2826 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=132460 $Y=49090 $D=28
M2115 2834 398 2832 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=132780 $Y=49090 $D=28
M2116 VSS 543 2834 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=133100 $Y=49090 $D=28
M2117 VSS clk 2825 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=134080 $Y=48840 $D=28
M2118 2828 2825 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=134590 $Y=48940 $D=28
M2119 2836 2828 2826 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=135610 $Y=49010 $D=28
M2120 2837 2827 2836 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=135930 $Y=49010 $D=28
M2121 VSS 543 2837 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=136250 $Y=49010 $D=28
M2122 2827 2826 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=136710 $Y=48870 $D=28
M2123 2829 2828 2827 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=137270 $Y=48870 $D=28
M2124 2839 2825 2829 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=137830 $Y=49110 $D=28
M2125 VSS 2831 2839 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=138150 $Y=49110 $D=28
M2126 2840 543 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=138590 $Y=49090 $D=28
M2127 2831 2829 2840 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=138910 $Y=49090 $D=28
M2128 2830 2831 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=139230 $Y=48390 $D=28
M2129 VSS 2830 930 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=140130 $Y=49070 $D=28
M2130 data_out[6] 2831 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=140630 $Y=49070 $D=28
M2131 2848 2841 2842 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=138460 $Y=53910 $D=28
M2132 2850 538 2848 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=138780 $Y=53910 $D=28
M2133 VSS 544 2850 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=139100 $Y=53910 $D=28
M2134 VSS clk 2841 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=140080 $Y=54060 $D=28
M2135 2844 2841 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=140590 $Y=54060 $D=28
M2136 2852 2844 2842 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=141610 $Y=53990 $D=28
M2137 2853 2843 2852 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=141930 $Y=53990 $D=28
M2138 VSS 544 2853 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=142250 $Y=53990 $D=28
M2139 2843 2842 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=142710 $Y=54130 $D=28
M2140 2845 2844 2843 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=143270 $Y=54130 $D=28
M2141 2855 2841 2845 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=143830 $Y=53890 $D=28
M2142 VSS 2847 2855 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=144150 $Y=53890 $D=28
M2143 2856 544 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=144590 $Y=53890 $D=28
M2144 2847 2845 2856 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=144910 $Y=53890 $D=28
M2145 2846 2847 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=145230 $Y=54610 $D=28
M2146 VSS 2846 931 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=146130 $Y=53890 $D=28
M2147 data_out[7] 2847 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=146630 $Y=53890 $D=28
M2148 2864 2857 2858 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=141260 $Y=46710 $D=28
M2149 2866 367 2864 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=141580 $Y=46710 $D=28
M2150 VSS 544 2866 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=141900 $Y=46710 $D=28
M2151 VSS clk 2857 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=142880 $Y=46860 $D=28
M2152 2860 2857 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=143390 $Y=46860 $D=28
M2153 2868 2860 2858 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=144410 $Y=46790 $D=28
M2154 2869 2859 2868 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=144730 $Y=46790 $D=28
M2155 VSS 544 2869 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=145050 $Y=46790 $D=28
M2156 2859 2858 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=145510 $Y=46930 $D=28
M2157 2861 2860 2859 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=146070 $Y=46930 $D=28
M2158 2871 2857 2861 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=146630 $Y=46690 $D=28
M2159 VSS 2863 2871 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=146950 $Y=46690 $D=28
M2160 2872 544 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=147390 $Y=46690 $D=28
M2161 2863 2861 2872 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=147710 $Y=46690 $D=28
M2162 2862 2863 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=148030 $Y=47410 $D=28
M2163 VSS 2862 932 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=148930 $Y=46690 $D=28
M2164 data_out[5] 2863 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=149430 $Y=46690 $D=28
M2165 2880 2873 2874 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=144060 $Y=20290 $D=28
M2166 2882 563 2880 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=144380 $Y=20290 $D=28
M2167 VSS 564 2882 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=144700 $Y=20290 $D=28
M2168 VSS clk 2873 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=145680 $Y=20040 $D=28
M2169 2876 2873 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=146190 $Y=20140 $D=28
M2170 2884 2876 2874 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=147210 $Y=20210 $D=28
M2171 2885 2875 2884 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=147530 $Y=20210 $D=28
M2172 VSS 564 2885 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=147850 $Y=20210 $D=28
M2173 2875 2874 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=148310 $Y=20070 $D=28
M2174 2877 2876 2875 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=148870 $Y=20070 $D=28
M2175 2887 2873 2877 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=149430 $Y=20310 $D=28
M2176 VSS 2879 2887 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=149750 $Y=20310 $D=28
M2177 2888 564 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=150190 $Y=20290 $D=28
M2178 2879 2877 2888 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=150510 $Y=20290 $D=28
M2179 2878 2879 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=150830 $Y=19590 $D=28
M2180 VSS 2878 933 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=151730 $Y=20270 $D=28
M2181 result[24] 2879 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=152230 $Y=20270 $D=28
M2182 2896 2889 2890 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=144060 $Y=39510 $D=28
M2183 2898 176 2896 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=144380 $Y=39510 $D=28
M2184 VSS 544 2898 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=144700 $Y=39510 $D=28
M2185 VSS clk 2889 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=145680 $Y=39660 $D=28
M2186 2892 2889 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=146190 $Y=39660 $D=28
M2187 2900 2892 2890 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=147210 $Y=39590 $D=28
M2188 2901 2891 2900 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=147530 $Y=39590 $D=28
M2189 VSS 544 2901 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=147850 $Y=39590 $D=28
M2190 2891 2890 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=148310 $Y=39730 $D=28
M2191 2893 2892 2891 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=148870 $Y=39730 $D=28
M2192 2903 2889 2893 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=149430 $Y=39490 $D=28
M2193 VSS 2895 2903 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=149750 $Y=39490 $D=28
M2194 2904 544 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=150190 $Y=39490 $D=28
M2195 2895 2893 2904 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=150510 $Y=39490 $D=28
M2196 2894 2895 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=150830 $Y=40210 $D=28
M2197 VSS 2894 934 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=151730 $Y=39490 $D=28
M2198 data_out[4] 2895 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=152230 $Y=39490 $D=28
M2199 2912 2905 2906 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=148060 $Y=25110 $D=28
M2200 2914 654 2912 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=148380 $Y=25110 $D=28
M2201 VSS 662 2914 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=148700 $Y=25110 $D=28
M2202 VSS clk 2905 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=149680 $Y=25260 $D=28
M2203 2908 2905 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=150190 $Y=25260 $D=28
M2204 2916 2908 2906 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=151210 $Y=25190 $D=28
M2205 2917 2907 2916 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=151530 $Y=25190 $D=28
M2206 VSS 662 2917 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=151850 $Y=25190 $D=28
M2207 2907 2906 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=152310 $Y=25330 $D=28
M2208 2909 2908 2907 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=152870 $Y=25330 $D=28
M2209 2919 2905 2909 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=153430 $Y=25090 $D=28
M2210 VSS 2911 2919 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=153750 $Y=25090 $D=28
M2211 2920 662 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=154190 $Y=25090 $D=28
M2212 2911 2909 2920 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=154510 $Y=25090 $D=28
M2213 2910 2911 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=154830 $Y=25810 $D=28
M2214 VSS 2910 935 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=155730 $Y=25090 $D=28
M2215 result[23] 2911 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=156230 $Y=25090 $D=28
M2216 2928 2921 2922 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=156060 $Y=10710 $D=28
M2217 2930 621 2928 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=156380 $Y=10710 $D=28
M2218 VSS 665 2930 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=156700 $Y=10710 $D=28
M2219 VSS clk 2921 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=157680 $Y=10860 $D=28
M2220 2924 2921 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=158190 $Y=10860 $D=28
M2221 2932 2924 2922 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=159210 $Y=10790 $D=28
M2222 2933 2923 2932 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=159530 $Y=10790 $D=28
M2223 VSS 665 2933 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=159850 $Y=10790 $D=28
M2224 2923 2922 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=160310 $Y=10930 $D=28
M2225 2925 2924 2923 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=160870 $Y=10930 $D=28
M2226 2935 2921 2925 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=161430 $Y=10690 $D=28
M2227 VSS 2927 2935 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=161750 $Y=10690 $D=28
M2228 2936 665 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=162190 $Y=10690 $D=28
M2229 2927 2925 2936 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=162510 $Y=10690 $D=28
M2230 2926 2927 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=162830 $Y=11410 $D=28
M2231 VSS 2926 936 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=163730 $Y=10690 $D=28
M2232 result[22] 2927 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=164230 $Y=10690 $D=28
M2233 2944 2937 2938 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=159660 $Y=20290 $D=28
M2234 2946 678 2944 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=159980 $Y=20290 $D=28
M2235 VSS 638 2946 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=160300 $Y=20290 $D=28
M2236 VSS clk 2937 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=161280 $Y=20040 $D=28
M2237 2940 2937 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=161790 $Y=20140 $D=28
M2238 2948 2940 2938 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=162810 $Y=20210 $D=28
M2239 2949 2939 2948 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=163130 $Y=20210 $D=28
M2240 VSS 638 2949 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=163450 $Y=20210 $D=28
M2241 2939 2938 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=163910 $Y=20070 $D=28
M2242 2941 2940 2939 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=164470 $Y=20070 $D=28
M2243 2951 2937 2941 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=165030 $Y=20310 $D=28
M2244 VSS 2943 2951 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=165350 $Y=20310 $D=28
M2245 2952 638 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=165790 $Y=20290 $D=28
M2246 2943 2941 2952 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=166110 $Y=20290 $D=28
M2247 2942 2943 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=166430 $Y=19590 $D=28
M2248 VSS 2942 937 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=167330 $Y=20270 $D=28
M2249 result[27] 2943 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=167830 $Y=20270 $D=28
M2250 2960 2953 2954 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=160860 $Y=13090 $D=28
M2251 2962 643 2960 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=161180 $Y=13090 $D=28
M2252 VSS 665 2962 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=161500 $Y=13090 $D=28
M2253 VSS clk 2953 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=162480 $Y=12840 $D=28
M2254 2956 2953 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=162990 $Y=12940 $D=28
M2255 2964 2956 2954 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=164010 $Y=13010 $D=28
M2256 2965 2955 2964 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=164330 $Y=13010 $D=28
M2257 VSS 665 2965 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=164650 $Y=13010 $D=28
M2258 2955 2954 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=165110 $Y=12870 $D=28
M2259 2957 2956 2955 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=165670 $Y=12870 $D=28
M2260 2967 2953 2957 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=166230 $Y=13110 $D=28
M2261 VSS 2959 2967 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=166550 $Y=13110 $D=28
M2262 2968 665 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=166990 $Y=13090 $D=28
M2263 2959 2957 2968 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=167310 $Y=13090 $D=28
M2264 2958 2959 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=167630 $Y=12390 $D=28
M2265 VSS 2958 938 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=168530 $Y=13070 $D=28
M2266 result[28] 2959 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=169030 $Y=13070 $D=28
M2267 2976 2969 2970 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=166460 $Y=10710 $D=28
M2268 2978 699 2976 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=166780 $Y=10710 $D=28
M2269 VSS 665 2978 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=167100 $Y=10710 $D=28
M2270 VSS clk 2969 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=168080 $Y=10860 $D=28
M2271 2972 2969 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=168590 $Y=10860 $D=28
M2272 2980 2972 2970 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=169610 $Y=10790 $D=28
M2273 2981 2971 2980 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=169930 $Y=10790 $D=28
M2274 VSS 665 2981 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=170250 $Y=10790 $D=28
M2275 2971 2970 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=170710 $Y=10930 $D=28
M2276 2973 2972 2971 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=171270 $Y=10930 $D=28
M2277 2983 2969 2973 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=171830 $Y=10690 $D=28
M2278 VSS 2975 2983 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=172150 $Y=10690 $D=28
M2279 2984 665 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=172590 $Y=10690 $D=28
M2280 2975 2973 2984 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=172910 $Y=10690 $D=28
M2281 2974 2975 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=173230 $Y=11410 $D=28
M2282 VSS 2974 939 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=174130 $Y=10690 $D=28
M2283 result[29] 2975 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=174630 $Y=10690 $D=28
M2284 2992 2985 2986 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=168060 $Y=17910 $D=28
M2285 2994 708 2992 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=168380 $Y=17910 $D=28
M2286 VSS 706 2994 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=168700 $Y=17910 $D=28
M2287 VSS clk 2985 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=169680 $Y=18060 $D=28
M2288 2988 2985 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=170190 $Y=18060 $D=28
M2289 2996 2988 2986 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=171210 $Y=17990 $D=28
M2290 2997 2987 2996 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=171530 $Y=17990 $D=28
M2291 VSS 706 2997 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=171850 $Y=17990 $D=28
M2292 2987 2986 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=172310 $Y=18130 $D=28
M2293 2989 2988 2987 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=172870 $Y=18130 $D=28
M2294 2999 2985 2989 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=173430 $Y=17890 $D=28
M2295 VSS 2991 2999 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=173750 $Y=17890 $D=28
M2296 3000 706 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=174190 $Y=17890 $D=28
M2297 2991 2989 3000 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=174510 $Y=17890 $D=28
M2298 2990 2991 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=174830 $Y=18610 $D=28
M2299 VSS 2990 940 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=175730 $Y=17890 $D=28
M2300 result[30] 2991 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=176230 $Y=17890 $D=28
M2301 3008 3001 3002 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=176060 $Y=10710 $D=28
M2302 3010 740 3008 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=176380 $Y=10710 $D=28
M2303 VSS 665 3010 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=176700 $Y=10710 $D=28
M2304 VSS clk 3001 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=177680 $Y=10860 $D=28
M2305 3004 3001 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=178190 $Y=10860 $D=28
M2306 3012 3004 3002 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=179210 $Y=10790 $D=28
M2307 3013 3003 3012 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=179530 $Y=10790 $D=28
M2308 VSS 665 3013 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=179850 $Y=10790 $D=28
M2309 3003 3002 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=180310 $Y=10930 $D=28
M2310 3005 3004 3003 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=180870 $Y=10930 $D=28
M2311 3015 3001 3005 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=181430 $Y=10690 $D=28
M2312 VSS 3007 3015 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=181750 $Y=10690 $D=28
M2313 3016 665 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=182190 $Y=10690 $D=28
M2314 3007 3005 3016 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=182510 $Y=10690 $D=28
M2315 3006 3007 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=182830 $Y=11410 $D=28
M2316 VSS 3006 941 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=183730 $Y=10690 $D=28
M2317 result[31] 3007 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=184230 $Y=10690 $D=28
M2318 VSS 80 3017 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=18040 $Y=68290 $D=28
M2319 3017 60 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=18520 $Y=68290 $D=28
M2320 802 50 3017 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=19000 $Y=68290 $D=28
M2321 VSS 220 3019 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=60440 $Y=55910 $D=28
M2322 3019 215 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=60920 $Y=55910 $D=28
M2323 229 210 3019 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=61400 $Y=55910 $D=28
M2324 VSS 412 3021 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=110040 $Y=53890 $D=28
M2325 3021 833 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=110520 $Y=53890 $D=28
M2326 835 414 3021 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=111000 $Y=53890 $D=28
M2327 VSS 417 3023 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=112040 $Y=63110 $D=28
M2328 3023 435 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=112520 $Y=63110 $D=28
M2329 420 476 3023 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=113000 $Y=63110 $D=28
M2330 VSS 458 3025 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=121640 $Y=34310 $D=28
M2331 3025 478 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=122120 $Y=34310 $D=28
M2332 459 477 3025 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=122600 $Y=34310 $D=28
M2333 VSS 492 3027 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=131240 $Y=39490 $D=28
M2334 3027 502 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=131720 $Y=39490 $D=28
M2335 506 517 3027 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=132200 $Y=39490 $D=28
M2336 VSS 522 3029 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=135240 $Y=32290 $D=28
M2337 3029 527 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=135720 $Y=32290 $D=28
M2338 546 551 3029 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=136200 $Y=32290 $D=28
M2339 VSS 528 3031 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=137240 $Y=32290 $D=28
M2340 3031 530 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=137720 $Y=32290 $D=28
M2341 537 536 3031 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=138200 $Y=32290 $D=28
M2342 VSS 600 3033 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=146040 $Y=48710 $D=28
M2343 3033 587 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=146520 $Y=48710 $D=28
M2344 606 580 3033 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=147000 $Y=48710 $D=28
M2345 VSS 581 3035 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=146440 $Y=55910 $D=28
M2346 3035 566 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=146920 $Y=55910 $D=28
M2347 559 607 3035 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=147400 $Y=55910 $D=28
M2348 VSS 591 3037 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=147240 $Y=34310 $D=28
M2349 3037 571 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=147720 $Y=34310 $D=28
M2350 596 585 3037 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=148200 $Y=34310 $D=28
M2351 VSS 626 3039 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=156040 $Y=61090 $D=28
M2352 3039 616 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=156520 $Y=61090 $D=28
M2353 687 627 3039 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=157000 $Y=61090 $D=28
M2354 VSS 783 3041 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=174840 $Y=61090 $D=28
M2355 3041 784 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=175320 $Y=61090 $D=28
M2356 775 736 3041 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=175800 $Y=61090 $D=28
M2357 VSS 703 3043 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.92e-13 pd=9.6e-07 ps=1.84e-06 nrd=0.3 nrs=0.533333 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=175640 $Y=48710 $D=28
M2358 3043 721 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=176120 $Y=48710 $D=28
M2359 727 724 3043 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=176600 $Y=48710 $D=28
M2360 22 70 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.728e-13 pd=1.6e-06 ps=1.68e-06 nrd=0.666667 nrs=0.75 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=17830 $Y=32290 $D=28
M2361 204 167 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.728e-13 pd=1.6e-06 ps=1.68e-06 nrd=0.666667 nrs=0.75 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=51030 $Y=17890 $D=28
M2362 286 285 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.728e-13 pd=1.6e-06 ps=1.68e-06 nrd=0.666667 nrs=0.75 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=75830 $Y=41630 $D=28
M2363 830 353 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.728e-13 pd=1.6e-06 ps=1.68e-06 nrd=0.666667 nrs=0.75 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=95430 $Y=70430 $D=28
M2364 584 850 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.728e-13 pd=1.6e-06 ps=1.68e-06 nrd=0.666667 nrs=0.75 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=139830 $Y=12830 $D=28
M2365 719 674 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.728e-13 pd=1.6e-06 ps=1.68e-06 nrd=0.666667 nrs=0.75 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=175430 $Y=70430 $D=28
M2366 112 89 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.24696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=27300 $Y=41190 $D=28
M2367 VSS 89 112 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.22525e-13 as=1.656e-13 pd=1.56208e-06 ps=1.28e-06 nrd=0.262908 nrs=0.195652 sa=8e-07 sb=7.66957e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=27780 $Y=41190 $D=28
M2368 112 89 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.7415e-13 pd=2.08e-06 ps=1.2225e-06 nrd=0.444444 nrs=0.335937 sa=1.36e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=28340 $Y=41390 $D=28
M2369 201 172 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.24696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=50900 $Y=75490 $D=28
M2370 VSS 172 201 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.22525e-13 as=1.656e-13 pd=1.56208e-06 ps=1.28e-06 nrd=0.262908 nrs=0.195652 sa=8e-07 sb=7.66957e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=51380 $Y=75490 $D=28
M2371 201 172 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.7415e-13 pd=2.08e-06 ps=1.2225e-06 nrd=0.444444 nrs=0.335937 sa=1.36e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=51940 $Y=75490 $D=28
M2372 263 201 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.24696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=60900 $Y=48390 $D=28
M2373 VSS 201 263 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.22525e-13 as=1.656e-13 pd=1.56208e-06 ps=1.28e-06 nrd=0.262908 nrs=0.195652 sa=8e-07 sb=7.66957e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=61380 $Y=48390 $D=28
M2374 263 201 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.7415e-13 pd=2.08e-06 ps=1.2225e-06 nrd=0.444444 nrs=0.335937 sa=1.36e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=61940 $Y=48590 $D=28
M2375 518 849 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.24696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=134100 $Y=62790 $D=28
M2376 VSS 849 518 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.22525e-13 as=1.656e-13 pd=1.56208e-06 ps=1.28e-06 nrd=0.262908 nrs=0.195652 sa=8e-07 sb=7.66957e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=134580 $Y=62790 $D=28
M2377 518 849 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.7415e-13 pd=2.08e-06 ps=1.2225e-06 nrd=0.444444 nrs=0.335937 sa=1.36e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=135140 $Y=62990 $D=28
M2378 562 849 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.24696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=135300 $Y=68290 $D=28
M2379 VSS 849 562 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.22525e-13 as=1.656e-13 pd=1.56208e-06 ps=1.28e-06 nrd=0.262908 nrs=0.195652 sa=8e-07 sb=7.66957e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=135780 $Y=68290 $D=28
M2380 562 849 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.7415e-13 pd=2.08e-06 ps=1.2225e-06 nrd=0.444444 nrs=0.335937 sa=1.36e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=136340 $Y=68290 $D=28
M2381 742 523 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.24696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=169300 $Y=33990 $D=28
M2382 VSS 523 742 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.22525e-13 as=1.656e-13 pd=1.56208e-06 ps=1.28e-06 nrd=0.262908 nrs=0.195652 sa=8e-07 sb=7.66957e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=169780 $Y=33990 $D=28
M2383 742 523 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.7415e-13 pd=2.08e-06 ps=1.2225e-06 nrd=0.444444 nrs=0.335937 sa=1.36e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=170340 $Y=34190 $D=28
M2384 729 523 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.24696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=173300 $Y=62790 $D=28
M2385 VSS 523 729 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.22525e-13 as=1.656e-13 pd=1.56208e-06 ps=1.28e-06 nrd=0.262908 nrs=0.195652 sa=8e-07 sb=7.66957e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=173780 $Y=62790 $D=28
M2386 729 523 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.7415e-13 pd=2.08e-06 ps=1.2225e-06 nrd=0.444444 nrs=0.335937 sa=1.36e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=174340 $Y=62990 $D=28
M2387 VSS 85 3045 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.952e-13 pd=1.32573e-06 ps=1.86e-06 nrd=0.47082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=25680 $Y=70300 $D=28
M2388 3045 81 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=8.8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=26240 $Y=70300 $D=28
M2389 VSS 81 3045 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.47082 nrs=0.295082 sa=1.36e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=26720 $Y=70300 $D=28
M2390 3045 85 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=1.92e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=27280 $Y=70300 $D=28
M2391 885 91 3045 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=27760 $Y=70300 $D=28
M2392 3045 91 885 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=28240 $Y=70300 $D=28
M2393 VSS 218 3048 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.952e-13 pd=1.32573e-06 ps=1.86e-06 nrd=0.47082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=58080 $Y=53890 $D=28
M2394 3048 221 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=8.8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=58640 $Y=53890 $D=28
M2395 VSS 221 3048 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.47082 nrs=0.295082 sa=1.36e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=59120 $Y=53890 $D=28
M2396 3048 218 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=1.92e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=59680 $Y=53890 $D=28
M2397 220 247 3048 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=60160 $Y=53890 $D=28
M2398 3048 247 220 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=60640 $Y=53890 $D=28
M2399 VSS 281 3051 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.952e-13 pd=1.32573e-06 ps=1.86e-06 nrd=0.47082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=62880 $Y=19900 $D=28
M2400 3051 249 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=8.8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=63440 $Y=19900 $D=28
M2401 VSS 249 3051 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.47082 nrs=0.295082 sa=1.36e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=63920 $Y=19900 $D=28
M2402 3051 281 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=1.92e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=64480 $Y=19900 $D=28
M2403 235 258 3051 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=64960 $Y=19900 $D=28
M2404 3051 258 235 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=65440 $Y=19900 $D=28
M2405 VSS 439 3054 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.952e-13 pd=1.32573e-06 ps=1.86e-06 nrd=0.47082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=116480 $Y=70300 $D=28
M2406 3054 435 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=8.8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=117040 $Y=70300 $D=28
M2407 VSS 435 3054 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.47082 nrs=0.295082 sa=1.36e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=117520 $Y=70300 $D=28
M2408 3054 439 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=1.92e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=118080 $Y=70300 $D=28
M2409 840 468 3054 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=118560 $Y=70300 $D=28
M2410 3054 468 840 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=119040 $Y=70300 $D=28
M2411 VSS 574 3057 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.952e-13 pd=1.32573e-06 ps=1.86e-06 nrd=0.47082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=157280 $Y=55900 $D=28
M2412 3057 637 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=8.8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=157840 $Y=55900 $D=28
M2413 VSS 637 3057 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.47082 nrs=0.295082 sa=1.36e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=158320 $Y=55900 $D=28
M2414 3057 574 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=1.92e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=158880 $Y=55900 $D=28
M2415 664 649 3057 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=159360 $Y=55900 $D=28
M2416 3057 649 664 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=159840 $Y=55900 $D=28
M2417 VSS 648 3060 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.952e-13 pd=1.32573e-06 ps=1.86e-06 nrd=0.47082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=158480 $Y=61090 $D=28
M2418 3060 659 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=8.8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=159040 $Y=61090 $D=28
M2419 VSS 659 3060 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.47082 nrs=0.295082 sa=1.36e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=159520 $Y=61090 $D=28
M2420 3060 648 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=1.92e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=160080 $Y=61090 $D=28
M2421 674 640 3060 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=160560 $Y=61090 $D=28
M2422 3060 640 674 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=161040 $Y=61090 $D=28
M2423 VSS 686 3063 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.952e-13 pd=1.32573e-06 ps=1.86e-06 nrd=0.47082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=170880 $Y=68290 $D=28
M2424 3063 719 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=8.8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=171440 $Y=68290 $D=28
M2425 VSS 719 3063 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.47082 nrs=0.295082 sa=1.36e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=171920 $Y=68290 $D=28
M2426 3063 686 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=1.92e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=172480 $Y=68290 $D=28
M2427 758 692 3063 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=172960 $Y=68290 $D=28
M2428 3063 692 758 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=173440 $Y=68290 $D=28
M2429 VSS 731 3066 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.952e-13 pd=1.32573e-06 ps=1.86e-06 nrd=0.47082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=172880 $Y=39490 $D=28
M2430 3066 690 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=8.8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=173440 $Y=39490 $D=28
M2431 VSS 690 3066 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.75192e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.47082 nrs=0.295082 sa=1.36e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=173920 $Y=39490 $D=28
M2432 3066 731 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.75192e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.47082 sa=1.92e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=174480 $Y=39490 $D=28
M2433 741 735 3066 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=174960 $Y=39490 $D=28
M2434 3066 735 741 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=175440 $Y=39490 $D=28
M2435 80 69 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=3.1188e-13 pd=1.28e-06 ps=2.37667e-06 nrd=0.195652 nrs=0.368478 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=22120 $Y=62790 $D=28
M2436 VSS 121 80 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8.4e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=22600 $Y=62790 $D=28
M2437 80 121 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.08475e-13 pd=1.28e-06 ps=1.41472e-06 nrd=0.195652 nrs=0.246308 sa=1.4e-06 sb=1.24e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=23160 $Y=62790 $D=28
M2438 VSS 69 80 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.15112e-13 as=1.656e-13 pd=1.97143e-06 ps=1.28e-06 nrd=0.490444 nrs=0.195652 sa=1.88e-06 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=23640 $Y=62790 $D=28
M2439 119 125 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=3.1188e-13 pd=1.28e-06 ps=2.37667e-06 nrd=0.195652 nrs=0.368478 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=35320 $Y=26790 $D=28
M2440 VSS 130 119 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8.4e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=35800 $Y=26790 $D=28
M2441 119 130 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.08475e-13 pd=1.28e-06 ps=1.41472e-06 nrd=0.195652 nrs=0.246308 sa=1.4e-06 sb=1.24e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=36360 $Y=26790 $D=28
M2442 VSS 125 119 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.15112e-13 as=1.656e-13 pd=1.97143e-06 ps=1.28e-06 nrd=0.490444 nrs=0.195652 sa=1.88e-06 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=36840 $Y=26790 $D=28
M2443 81 191 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=3.1188e-13 pd=1.28e-06 ps=2.37667e-06 nrd=0.195652 nrs=0.368478 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=36920 $Y=75490 $D=28
M2444 VSS 238 81 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8.4e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=37400 $Y=75490 $D=28
M2445 81 238 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.08475e-13 pd=1.28e-06 ps=1.41472e-06 nrd=0.195652 nrs=0.246308 sa=1.4e-06 sb=1.24e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=37960 $Y=75490 $D=28
M2446 VSS 191 81 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.15112e-13 as=1.656e-13 pd=1.97143e-06 ps=1.28e-06 nrd=0.490444 nrs=0.195652 sa=1.88e-06 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=38440 $Y=75490 $D=28
M2447 366 308 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=3.1188e-13 pd=1.28e-06 ps=2.37667e-06 nrd=0.195652 nrs=0.368478 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=82120 $Y=75490 $D=28
M2448 VSS 347 366 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8.4e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=82600 $Y=75490 $D=28
M2449 366 347 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.08475e-13 pd=1.28e-06 ps=1.41472e-06 nrd=0.195652 nrs=0.246308 sa=1.4e-06 sb=1.24e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=83160 $Y=75490 $D=28
M2450 VSS 308 366 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.15112e-13 as=1.656e-13 pd=1.97143e-06 ps=1.28e-06 nrd=0.490444 nrs=0.195652 sa=1.88e-06 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=83640 $Y=75490 $D=28
M2451 473 353 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=3.1188e-13 pd=1.28e-06 ps=2.37667e-06 nrd=0.195652 nrs=0.368478 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=92520 $Y=75490 $D=28
M2452 VSS 366 473 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8.4e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=93000 $Y=75490 $D=28
M2453 473 366 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.08475e-13 pd=1.28e-06 ps=1.41472e-06 nrd=0.195652 nrs=0.246308 sa=1.4e-06 sb=1.24e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=93560 $Y=75490 $D=28
M2454 VSS 353 473 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.15112e-13 as=1.656e-13 pd=1.97143e-06 ps=1.28e-06 nrd=0.490444 nrs=0.195652 sa=1.88e-06 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=94040 $Y=75490 $D=28
M2455 490 846 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=3.1188e-13 pd=1.28e-06 ps=2.37667e-06 nrd=0.195652 nrs=0.368478 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=126920 $Y=69990 $D=28
M2456 VSS 417 490 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8.4e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=127400 $Y=69990 $D=28
M2457 490 417 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.08475e-13 pd=1.28e-06 ps=1.41472e-06 nrd=0.195652 nrs=0.246308 sa=1.4e-06 sb=1.24e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=127960 $Y=69990 $D=28
M2458 VSS 846 490 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.15112e-13 as=1.656e-13 pd=1.97143e-06 ps=1.28e-06 nrd=0.490444 nrs=0.195652 sa=1.88e-06 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=128440 $Y=69990 $D=28
M2459 508 485 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=3.1188e-13 pd=1.28e-06 ps=2.37667e-06 nrd=0.195652 nrs=0.368478 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=130120 $Y=55590 $D=28
M2460 VSS 521 508 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8.4e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=130600 $Y=55590 $D=28
M2461 508 521 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.08475e-13 pd=1.28e-06 ps=1.41472e-06 nrd=0.195652 nrs=0.246308 sa=1.4e-06 sb=1.24e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=131160 $Y=55590 $D=28
M2462 VSS 485 508 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.15112e-13 as=1.656e-13 pd=1.97143e-06 ps=1.28e-06 nrd=0.490444 nrs=0.195652 sa=1.88e-06 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=131640 $Y=55590 $D=28
M2463 694 681 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=3.1188e-13 pd=1.28e-06 ps=2.37667e-06 nrd=0.195652 nrs=0.368478 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=168520 $Y=41190 $D=28
M2464 VSS 700 694 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8.4e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=169000 $Y=41190 $D=28
M2465 694 700 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.08475e-13 pd=1.28e-06 ps=1.41472e-06 nrd=0.195652 nrs=0.246308 sa=1.4e-06 sb=1.24e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=169560 $Y=41190 $D=28
M2466 VSS 681 694 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.15112e-13 as=1.656e-13 pd=1.97143e-06 ps=1.28e-06 nrd=0.490444 nrs=0.195652 sa=1.88e-06 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=170040 $Y=41190 $D=28
M2467 704 693 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=3.1188e-13 pd=1.28e-06 ps=2.37667e-06 nrd=0.195652 nrs=0.368478 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=172120 $Y=25090 $D=28
M2468 VSS 743 704 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8.4e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=172600 $Y=25090 $D=28
M2469 704 743 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.08475e-13 pd=1.28e-06 ps=1.41472e-06 nrd=0.195652 nrs=0.246308 sa=1.4e-06 sb=1.24e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=173160 $Y=25090 $D=28
M2470 VSS 693 704 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.15112e-13 as=1.656e-13 pd=1.97143e-06 ps=1.28e-06 nrd=0.490444 nrs=0.195652 sa=1.88e-06 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=173640 $Y=25090 $D=28
M2471 556 581 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.12e-14 as=1.27754e-13 pd=7.4e-07 ps=1.18154e-06 nrd=1.0625 nrs=2.21795 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=3.6e-15 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=142070 $Y=61360 $D=28
M2472 VSS 557 556 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.592e-13 as=6.12e-14 pd=1.72e-06 ps=7.4e-07 nrd=2.76389 nrs=1.0625 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=3.6e-15 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=142630 $Y=61360 $D=28
M2473 653 666 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.12e-14 as=1.27754e-13 pd=7.4e-07 ps=1.18154e-06 nrd=1.0625 nrs=2.21795 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=3.6e-15 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=164070 $Y=56000 $D=28
M2474 VSS 667 653 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.592e-13 as=6.12e-14 pd=1.72e-06 ps=7.4e-07 nrd=2.76389 nrs=1.0625 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=3.6e-15 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=164630 $Y=56000 $D=28
M2475 691 713 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.12e-14 as=1.27754e-13 pd=7.4e-07 ps=1.18154e-06 nrd=1.0625 nrs=2.21795 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=3.6e-15 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=165670 $Y=56000 $D=28
M2476 VSS 667 691 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.592e-13 as=6.12e-14 pd=1.72e-06 ps=7.4e-07 nrd=2.76389 nrs=1.0625 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=3.6e-15 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=166230 $Y=56000 $D=28
M2477 731 683 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.12e-14 as=1.27754e-13 pd=7.4e-07 ps=1.18154e-06 nrd=1.0625 nrs=2.21795 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=3.6e-15 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=171670 $Y=34400 $D=28
M2478 VSS 709 731 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.592e-13 as=6.12e-14 pd=1.72e-06 ps=7.4e-07 nrd=2.76389 nrs=1.0625 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=3.6e-15 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=172230 $Y=34400 $D=28
M2479 3101 14 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=3.123e-13 pd=8e-07 ps=2.52e-06 nrd=0.166667 nrs=0.8675 sa=3.9e-07 sb=1.06933e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=15290 $Y=53890 $D=28
M2480 45 13 3101 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29509e-13 as=6e-14 pd=1.13208e-06 ps=8e-07 nrd=0.359748 nrs=0.166667 sa=7.1e-07 sb=7.49333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=15610 $Y=53890 $D=28
M2481 VSS 38 45 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.748e-13 as=9.92906e-14 pd=2.42e-06 ps=8.67925e-07 nrd=1.29868 nrs=0.469237 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=16130 $Y=53890 $D=28
M2482 3103 443 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=3.123e-13 pd=8e-07 ps=2.52e-06 nrd=0.166667 nrs=0.8675 sa=3.9e-07 sb=1.06933e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=123690 $Y=68290 $D=28
M2483 468 465 3103 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29509e-13 as=6e-14 pd=1.13208e-06 ps=8e-07 nrd=0.359748 nrs=0.166667 sa=7.1e-07 sb=7.49333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=124010 $Y=68290 $D=28
M2484 VSS 467 468 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.748e-13 as=9.92906e-14 pd=2.42e-06 ps=8.67925e-07 nrd=1.29868 nrs=0.469237 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=124530 $Y=68290 $D=28
M2485 3105 484 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=3.123e-13 pd=8e-07 ps=2.52e-06 nrd=0.166667 nrs=0.8675 sa=3.9e-07 sb=1.06933e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=128890 $Y=32290 $D=28
M2486 527 501 3105 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29509e-13 as=6e-14 pd=1.13208e-06 ps=8e-07 nrd=0.359748 nrs=0.166667 sa=7.1e-07 sb=7.49333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=129210 $Y=32290 $D=28
M2487 VSS 847 527 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.748e-13 as=9.92906e-14 pd=2.42e-06 ps=8.67925e-07 nrd=1.29868 nrs=0.469237 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=129730 $Y=32290 $D=28
M2488 3107 515 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=3.123e-13 pd=8e-07 ps=2.52e-06 nrd=0.166667 nrs=0.8675 sa=3.9e-07 sb=1.06933e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=128890 $Y=34310 $D=28
M2489 530 506 3107 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29509e-13 as=6e-14 pd=1.13208e-06 ps=8e-07 nrd=0.359748 nrs=0.166667 sa=7.1e-07 sb=7.49333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=129210 $Y=34310 $D=28
M2490 VSS 851 530 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.748e-13 as=9.92906e-14 pd=2.42e-06 ps=8.67925e-07 nrd=1.29868 nrs=0.469237 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=129730 $Y=34450 $D=28
M2491 3109 914 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=3.123e-13 pd=8e-07 ps=2.52e-06 nrd=0.166667 nrs=0.8675 sa=3.9e-07 sb=1.06933e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=140490 $Y=32290 $D=28
M2492 551 558 3109 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29509e-13 as=6e-14 pd=1.13208e-06 ps=8e-07 nrd=0.359748 nrs=0.166667 sa=7.1e-07 sb=7.49333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=140810 $Y=32290 $D=28
M2493 VSS 550 551 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.748e-13 as=9.92906e-14 pd=2.42e-06 ps=8.67925e-07 nrd=1.29868 nrs=0.469237 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=141330 $Y=32290 $D=28
M2494 3111 601 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=3.123e-13 pd=8e-07 ps=2.52e-06 nrd=0.166667 nrs=0.8675 sa=3.9e-07 sb=1.06933e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=150490 $Y=53890 $D=28
M2495 566 598 3111 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29509e-13 as=6e-14 pd=1.13208e-06 ps=8e-07 nrd=0.359748 nrs=0.166667 sa=7.1e-07 sb=7.49333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=150810 $Y=53890 $D=28
M2496 VSS 619 566 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.748e-13 as=9.92906e-14 pd=2.42e-06 ps=8.67925e-07 nrd=1.29868 nrs=0.469237 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=151330 $Y=53890 $D=28
M2497 3113 599 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=3.123e-13 pd=8e-07 ps=2.52e-06 nrd=0.166667 nrs=0.8675 sa=3.9e-07 sb=1.06933e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=151290 $Y=61090 $D=28
M2498 627 602 3113 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29509e-13 as=6e-14 pd=1.13208e-06 ps=8e-07 nrd=0.359748 nrs=0.166667 sa=7.1e-07 sb=7.49333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=151610 $Y=61090 $D=28
M2499 VSS 603 627 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.748e-13 as=9.92906e-14 pd=2.42e-06 ps=8.67925e-07 nrd=1.29868 nrs=0.469237 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=152130 $Y=61090 $D=28
M2500 3115 635 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=3.123e-13 pd=8e-07 ps=2.52e-06 nrd=0.166667 nrs=0.8675 sa=3.9e-07 sb=1.06933e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=154090 $Y=55910 $D=28
M2501 616 625 3115 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29509e-13 as=6e-14 pd=1.13208e-06 ps=8e-07 nrd=0.359748 nrs=0.166667 sa=7.1e-07 sb=7.49333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=154410 $Y=55910 $D=28
M2502 VSS 629 616 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.748e-13 as=9.92906e-14 pd=2.42e-06 ps=8.67925e-07 nrd=1.29868 nrs=0.469237 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=154930 $Y=56050 $D=28
M2503 3117 685 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=3.123e-13 pd=8e-07 ps=2.52e-06 nrd=0.166667 nrs=0.8675 sa=3.9e-07 sb=1.06933e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=168890 $Y=55910 $D=28
M2504 721 687 3117 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29509e-13 as=6e-14 pd=1.13208e-06 ps=8e-07 nrd=0.359748 nrs=0.166667 sa=7.1e-07 sb=7.49333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=169210 $Y=55910 $D=28
M2505 VSS 718 721 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.748e-13 as=9.92906e-14 pd=2.42e-06 ps=8.67925e-07 nrd=1.29868 nrs=0.469237 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=169730 $Y=56050 $D=28
M2506 3119 862 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=3.123e-13 pd=8e-07 ps=2.52e-06 nrd=0.166667 nrs=0.8675 sa=3.9e-07 sb=1.06933e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=170890 $Y=55910 $D=28
M2507 725 684 3119 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29509e-13 as=6e-14 pd=1.13208e-06 ps=8e-07 nrd=0.359748 nrs=0.166667 sa=7.1e-07 sb=7.49333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=171210 $Y=55910 $D=28
M2508 VSS 698 725 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.748e-13 as=9.92906e-14 pd=2.42e-06 ps=8.67925e-07 nrd=1.29868 nrs=0.469237 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=171730 $Y=56050 $D=28
M2509 3121 773 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=3.123e-13 pd=8e-07 ps=2.52e-06 nrd=0.166667 nrs=0.8675 sa=3.9e-07 sb=1.06933e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=171290 $Y=61090 $D=28
M2510 714 732 3121 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29509e-13 as=6e-14 pd=1.13208e-06 ps=8e-07 nrd=0.359748 nrs=0.166667 sa=7.1e-07 sb=7.49333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=171610 $Y=61090 $D=28
M2511 VSS 747 714 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.748e-13 as=9.92906e-14 pd=2.42e-06 ps=8.67925e-07 nrd=1.29868 nrs=0.469237 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=172130 $Y=61090 $D=28
M2512 VSS weight_in[1] 3122 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66817e-13 as=2.856e-13 pd=1.17915e-06 ps=2.2e-06 nrd=0.360763 nrs=0.617647 sa=4.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=25720 $Y=75490 $D=28
M2513 86 3122 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.25694e-13 pd=1.28e-06 ps=1.59532e-06 nrd=0.195652 nrs=0.266651 sa=8.18261e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=26280 $Y=75490 $D=28
M2514 VSS 3122 86 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.29826e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=26760 $Y=75490 $D=28
M2515 VSS 101 3123 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66817e-13 as=2.856e-13 pd=1.17915e-06 ps=2.2e-06 nrd=0.360763 nrs=0.617647 sa=4.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=29320 $Y=27030 $D=28
M2516 129 3123 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.25694e-13 pd=1.28e-06 ps=1.59532e-06 nrd=0.195652 nrs=0.266651 sa=8.18261e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=29880 $Y=26790 $D=28
M2517 VSS 3123 129 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.29826e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=30360 $Y=26790 $D=28
M2518 VSS 127 3124 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66817e-13 as=2.856e-13 pd=1.17915e-06 ps=2.2e-06 nrd=0.360763 nrs=0.617647 sa=4.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=30920 $Y=34230 $D=28
M2519 192 3124 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.25694e-13 pd=1.28e-06 ps=1.59532e-06 nrd=0.195652 nrs=0.266651 sa=8.18261e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=31480 $Y=33990 $D=28
M2520 VSS 3124 192 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.29826e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=31960 $Y=33990 $D=28
M2521 VSS 98 3125 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66817e-13 as=2.856e-13 pd=1.17915e-06 ps=2.2e-06 nrd=0.360763 nrs=0.617647 sa=4.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=37720 $Y=61090 $D=28
M2522 151 3125 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.25694e-13 pd=1.28e-06 ps=1.59532e-06 nrd=0.195652 nrs=0.266651 sa=8.18261e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=38280 $Y=61090 $D=28
M2523 VSS 3125 151 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.29826e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=38760 $Y=61090 $D=28
M2524 VSS 187 3126 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66817e-13 as=2.856e-13 pd=1.17915e-06 ps=2.2e-06 nrd=0.360763 nrs=0.617647 sa=4.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=69720 $Y=46690 $D=28
M2525 283 3126 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.25694e-13 pd=1.28e-06 ps=1.59532e-06 nrd=0.195652 nrs=0.266651 sa=8.18261e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=70280 $Y=46690 $D=28
M2526 VSS 3126 283 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.29826e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=70760 $Y=46690 $D=28
M2527 VSS 263 3127 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66817e-13 as=2.856e-13 pd=1.17915e-06 ps=2.2e-06 nrd=0.360763 nrs=0.617647 sa=4.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=70520 $Y=34230 $D=28
M2528 170 3127 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.25694e-13 pd=1.28e-06 ps=1.59532e-06 nrd=0.195652 nrs=0.266651 sa=8.18261e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=71080 $Y=33990 $D=28
M2529 VSS 3127 170 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.29826e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=71560 $Y=33990 $D=28
M2530 VSS 263 3128 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66817e-13 as=2.856e-13 pd=1.17915e-06 ps=2.2e-06 nrd=0.360763 nrs=0.617647 sa=4.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=72520 $Y=46690 $D=28
M2531 307 3128 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.25694e-13 pd=1.28e-06 ps=1.59532e-06 nrd=0.195652 nrs=0.266651 sa=8.18261e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=73080 $Y=46690 $D=28
M2532 VSS 3128 307 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.29826e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=73560 $Y=46690 $D=28
M2533 VSS 171 3129 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66817e-13 as=2.856e-13 pd=1.17915e-06 ps=2.2e-06 nrd=0.360763 nrs=0.617647 sa=4.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=102520 $Y=48630 $D=28
M2534 398 3129 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.25694e-13 pd=1.28e-06 ps=1.59532e-06 nrd=0.195652 nrs=0.266651 sa=8.18261e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=103080 $Y=48390 $D=28
M2535 VSS 3129 398 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.29826e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=103560 $Y=48390 $D=28
M2536 VSS 584 3130 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66817e-13 as=2.856e-13 pd=1.17915e-06 ps=2.2e-06 nrd=0.360763 nrs=0.617647 sa=4.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=148120 $Y=17890 $D=28
M2537 638 3130 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.25694e-13 pd=1.28e-06 ps=1.59532e-06 nrd=0.195652 nrs=0.266651 sa=8.18261e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=148680 $Y=17890 $D=28
M2538 VSS 3130 638 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.29826e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=149160 $Y=17890 $D=28
M2539 VSS 641 3131 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.66817e-13 as=2.856e-13 pd=1.17915e-06 ps=2.2e-06 nrd=0.360763 nrs=0.617647 sa=4.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=170520 $Y=32290 $D=28
M2540 706 3131 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.25694e-13 pd=1.28e-06 ps=1.59532e-06 nrd=0.195652 nrs=0.266651 sa=8.18261e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=171080 $Y=32290 $D=28
M2541 VSS 3131 706 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.656e-13 pd=2.37667e-06 ps=1.28e-06 nrd=0.368478 nrs=0.195652 sa=1.29826e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=171560 $Y=32290 $D=28
M2542 VSS 11 3132 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=8860 $Y=32290 $D=28
M2543 23 3132 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=9440 $Y=32290 $D=28
M2544 VSS data_in[4] 3133 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=8860 $Y=49110 $D=28
M2545 136 3133 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=9440 $Y=48830 $D=28
M2546 VSS data_in[6] 3134 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=8860 $Y=61090 $D=28
M2547 797 3134 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=9440 $Y=61090 $D=28
M2548 VSS data_in[3] 3135 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=10860 $Y=34710 $D=28
M2549 127 3135 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=11440 $Y=34430 $D=28
M2550 VSS 85 3136 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=13260 $Y=68290 $D=28
M2551 50 3136 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=13840 $Y=68290 $D=28
M2552 VSS rst_n 3137 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=19260 $Y=75490 $D=28
M2553 32 3137 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=19840 $Y=75490 $D=28
M2554 VSS 803 3138 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=23260 $Y=70710 $D=28
M2555 58 3138 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=23840 $Y=70430 $D=28
M2556 VSS 131 3139 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=46460 $Y=49110 $D=28
M2557 180 3139 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=47040 $Y=48830 $D=28
M2558 VSS 128 3140 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=48460 $Y=10690 $D=28
M2559 202 3140 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=49040 $Y=10690 $D=28
M2560 VSS 129 3141 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=58460 $Y=25090 $D=28
M2561 217 3141 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=59040 $Y=25090 $D=28
M2562 VSS 271 3142 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=61260 $Y=20310 $D=28
M2563 11 3142 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=61840 $Y=20030 $D=28
M2564 VSS 187 3143 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=63260 $Y=49110 $D=28
M2565 241 3143 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=63840 $Y=48830 $D=28
M2566 VSS 202 3144 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=64860 $Y=13110 $D=28
M2567 252 3144 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=65440 $Y=12830 $D=28
M2568 VSS 256 3145 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=71660 $Y=20310 $D=28
M2569 271 3145 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=72240 $Y=20030 $D=28
M2570 VSS 49 3146 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=73660 $Y=25090 $D=28
M2571 287 3146 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=74240 $Y=25090 $D=28
M2572 VSS 318 3147 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=82460 $Y=20310 $D=28
M2573 256 3147 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=83040 $Y=20030 $D=28
M2574 VSS 303 3148 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=85660 $Y=32290 $D=28
M2575 329 3148 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=86240 $Y=32290 $D=28
M2576 VSS 186 3149 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=86860 $Y=53890 $D=28
M2577 538 3149 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=87440 $Y=53890 $D=28
M2578 VSS 358 3150 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=97660 $Y=63510 $D=28
M2579 376 3150 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=98240 $Y=63230 $D=28
M2580 VSS 399 3151 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=105260 $Y=17890 $D=28
M2581 389 3151 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=105840 $Y=17890 $D=28
M2582 VSS 407 3152 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=106460 $Y=32290 $D=28
M2583 425 3152 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=107040 $Y=32290 $D=28
M2584 VSS 407 3153 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=108060 $Y=25090 $D=28
M2585 374 3153 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=108640 $Y=25090 $D=28
M2586 VSS 409 3154 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=108460 $Y=53890 $D=28
M2587 437 3154 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=109040 $Y=53890 $D=28
M2588 VSS 437 3155 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=117660 $Y=56310 $D=28
M2589 485 3155 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=118240 $Y=56030 $D=28
M2590 VSS 396 3156 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=121660 $Y=17890 $D=28
M2591 526 3156 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=122240 $Y=17890 $D=28
M2592 VSS 425 3157 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=124860 $Y=56310 $D=28
M2593 543 3157 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=125440 $Y=56030 $D=28
M2594 VSS 526 3158 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=135260 $Y=13110 $D=28
M2595 570 3158 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=135840 $Y=12830 $D=28
M2596 VSS 500 3159 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=141660 $Y=17890 $D=28
M2597 611 3159 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=142240 $Y=17890 $D=28
M2598 VSS 611 3160 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=147660 $Y=27510 $D=28
M2599 582 3160 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=148240 $Y=27230 $D=28
M2600 VSS 697 3161 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=152460 $Y=53890 $D=28
M2601 610 3161 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=153040 $Y=53890 $D=28
M2602 VSS 611 3162 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=153260 $Y=17890 $D=28
M2603 593 3162 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=153840 $Y=17890 $D=28
M2604 VSS 638 3163 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=159260 $Y=13110 $D=28
M2605 665 3163 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=159840 $Y=12830 $D=28
M2606 VSS 645 3164 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=161660 $Y=17890 $D=28
M2607 701 3164 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=162240 $Y=17890 $D=28
M2608 VSS 682 3165 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=169260 $Y=25090 $D=28
M2609 688 3165 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=169840 $Y=25090 $D=28
M2610 VSS data_in[1] 3166 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=8820 $Y=27150 $D=28
M2611 49 3166 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=9380 $Y=27020 $D=28
M2612 VSS 3166 49 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=9860 $Y=27020 $D=28
M2613 VSS 797 3167 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=8820 $Y=55950 $D=28
M2614 171 3167 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=9380 $Y=55820 $D=28
M2615 VSS 3167 171 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=9860 $Y=55820 $D=28
M2616 VSS 32 3168 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=20020 $Y=55950 $D=28
M2617 68 3168 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=20580 $Y=55820 $D=28
M2618 VSS 3168 68 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=21060 $Y=55820 $D=28
M2619 VSS weight_in[0] 3169 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=22420 $Y=75490 $D=28
M2620 97 3169 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=22980 $Y=75490 $D=28
M2621 VSS 3169 97 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=23460 $Y=75490 $D=28
M2622 VSS 82 3170 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=23620 $Y=34350 $D=28
M2623 74 3170 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=24180 $Y=34220 $D=28
M2624 VSS 3170 74 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=24660 $Y=34220 $D=28
M2625 VSS weight_in[2] 3171 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=28020 $Y=75490 $D=28
M2626 79 3171 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=28580 $Y=75490 $D=28
M2627 VSS 3171 79 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=29060 $Y=75490 $D=28
M2628 VSS 73 3172 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=30420 $Y=61090 $D=28
M2629 189 3172 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=30980 $Y=61090 $D=28
M2630 VSS 3172 189 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=31460 $Y=61090 $D=28
M2631 VSS 211 3173 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=36820 $Y=63150 $D=28
M2632 139 3173 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=37380 $Y=63020 $D=28
M2633 VSS 3173 139 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=37860 $Y=63020 $D=28
M2634 VSS weight_in[4] 3174 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=36820 $Y=70350 $D=28
M2635 153 3174 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=37380 $Y=70220 $D=28
M2636 VSS 3174 153 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=37860 $Y=70220 $D=28
M2637 VSS weight_in[5] 3175 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=44420 $Y=75490 $D=28
M2638 172 3175 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=44980 $Y=75490 $D=28
M2639 VSS 3175 172 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=45460 $Y=75490 $D=28
M2640 VSS weight_in[7] 3176 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=48820 $Y=75490 $D=28
M2641 187 3176 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=49380 $Y=75490 $D=28
M2642 VSS 3176 187 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=49860 $Y=75490 $D=28
M2643 VSS 141 3177 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=53620 $Y=32290 $D=28
M2644 254 3177 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=54180 $Y=32290 $D=28
M2645 VSS 3177 254 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=54660 $Y=32290 $D=28
M2646 VSS 213 3178 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=56020 $Y=53890 $D=28
M2647 218 3178 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=56580 $Y=53890 $D=28
M2648 VSS 3178 218 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=57060 $Y=53890 $D=28
M2649 VSS fire_in 3179 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=57620 $Y=75490 $D=28
M2650 306 3179 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=58180 $Y=75490 $D=28
M2651 VSS 3179 306 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=58660 $Y=75490 $D=28
M2652 VSS 187 3180 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=65220 $Y=41550 $D=28
M2653 240 3180 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=65780 $Y=41420 $D=28
M2654 VSS 3180 240 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=66260 $Y=41420 $D=28
M2655 VSS 252 3181 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=68020 $Y=12750 $D=28
M2656 299 3181 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=68580 $Y=12620 $D=28
M2657 VSS 3181 299 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=69060 $Y=12620 $D=28
M2658 VSS 246 3182 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=78420 $Y=55950 $D=28
M2659 295 3182 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=78980 $Y=55820 $D=28
M2660 VSS 3182 295 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=79460 $Y=55820 $D=28
M2661 VSS 157 3183 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=93620 $Y=39490 $D=28
M2662 367 3183 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=94180 $Y=39490 $D=28
M2663 VSS 3183 367 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=94660 $Y=39490 $D=28
M2664 VSS 348 3184 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=94820 $Y=55950 $D=28
M2665 360 3184 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=95380 $Y=55820 $D=28
M2666 VSS 3184 360 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=95860 $Y=55820 $D=28
M2667 VSS 371 3185 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=114820 $Y=10690 $D=28
M2668 428 3185 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=115380 $Y=10690 $D=28
M2669 VSS 3185 428 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=115860 $Y=10690 $D=28
M2670 VSS 408 3186 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=123220 $Y=17890 $D=28
M2671 491 3186 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=123780 $Y=17890 $D=28
M2672 VSS 3186 491 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=124260 $Y=17890 $D=28
M2673 VSS 428 3187 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=125220 $Y=17890 $D=28
M2674 479 3187 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=125780 $Y=17890 $D=28
M2675 VSS 3187 479 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=126260 $Y=17890 $D=28
M2676 VSS 491 3188 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=129220 $Y=12750 $D=28
M2677 500 3188 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=129780 $Y=12620 $D=28
M2678 VSS 3188 500 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=130260 $Y=12620 $D=28
M2679 VSS 638 3189 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=164420 $Y=25090 $D=28
M2680 662 3189 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=164980 $Y=25090 $D=28
M2681 VSS 3189 662 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=165460 $Y=25090 $D=28
M2682 VSS 689 3190 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.29606e-13 as=1.792e-13 pd=1.01248e-06 ps=1.76e-06 nrd=0.413286 nrs=0.571429 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=167620 $Y=27150 $D=28
M2683 693 3190 VSS VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.242e-13 as=1.59694e-13 pd=1.05e-06 ps=1.24752e-06 nrd=0.26087 nrs=0.33542 sa=7.76377e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=168180 $Y=27020 $D=28
M2684 VSS 3190 693 VSS lpnfet w=6.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.277e-13 as=1.242e-13 pd=2.04e-06 ps=1.05e-06 nrd=0.478261 nrs=0.26087 sa=1.25638e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=168660 $Y=27020 $D=28
M2685 27 26 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=16120 $Y=26790 $D=28
M2686 47 62 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=17320 $Y=26790 $D=28
M2687 76 117 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=23320 $Y=12390 $D=28
M2688 117 68 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=24520 $Y=12390 $D=28
M2689 303 302 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=78920 $Y=19590 $D=28
M2690 302 299 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=80120 $Y=19590 $D=28
M2691 344 316 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=93720 $Y=12390 $D=28
M2692 356 344 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=94920 $Y=12390 $D=28
M2693 525 492 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=134520 $Y=41190 $D=28
M2694 912 517 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=135720 $Y=41190 $D=28
M2695 534 502 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=136920 $Y=55590 $D=28
M2696 586 485 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=138120 $Y=55590 $D=28
M2697 655 620 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=157320 $Y=19590 $D=28
M2698 645 655 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=158520 $Y=19590 $D=28
M2699 658 662 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=159320 $Y=32290 $D=28
M2700 641 658 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=160520 $Y=32290 $D=28
M2701 667 669 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=163320 $Y=48390 $D=28
M2702 659 598 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=164520 $Y=48390 $D=28
M2703 860 688 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=166920 $Y=32290 $D=28
M2704 681 860 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=3.1188e-13 pd=2.48e-06 ps=2.37667e-06 nrd=0.347826 nrs=0.368478 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=168120 $Y=32290 $D=28
M2705 VSS clk 3191 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.624e-13 as=1.792e-13 pd=1.28121e-06 ps=1.76e-06 nrd=0.517857 nrs=0.571429 sa=3.2e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=119210 $Y=48630 $D=28
M2706 3195 clk VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=1.392e-13 pd=1.68e-06 ps=1.09818e-06 nrd=0.75 nrs=0.604167 sa=8.8e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=119770 $Y=48710 $D=28
M2707 VSS 508 3192 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37856e-13 as=1.536e-13 pd=1.0432e-06 ps=1.6e-06 nrd=0.598333 nrs=0.666667 sa=3.2e-07 sb=1.10333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=120900 $Y=48830 $D=28
M2708 3196 3191 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.12528e-13 pd=2.6e-06 ps=1.60827e-06 nrd=0.588751 nrs=0.388108 sa=6.97297e-07 sb=4.35676e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=121460 $Y=48570 $D=28
M2709 3201 3195 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7e-14 as=2.88e-13 pd=9e-07 ps=2.54e-06 nrd=0.142857 nrs=0.587755 sa=3.27429e-07 sb=1.36e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=122640 $Y=48710 $D=28
M2710 3193 3192 3201 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=7e-14 pd=1.06e-06 ps=9e-07 nrd=0.257143 nrs=0.142857 sa=6.47429e-07 sb=1.04e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=122960 $Y=48710 $D=28
M2711 3203 3192 3193 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7e-14 as=1.26e-13 pd=9e-07 ps=1.06e-06 nrd=0.142857 nrs=0.257143 sa=1.12743e-06 sb=5.6e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=123440 $Y=48710 $D=28
M2712 VSS 3195 3203 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.32857e-13 as=7e-14 pd=2.35714e-06 ps=9e-07 nrd=0.475219 nrs=0.142857 sa=1.44743e-06 sb=2.4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=123760 $Y=48710 $D=28
M2713 3205 3196 3193 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=8.4e-15 panw7=1.56e-14 panw8=0 panw9=0 panw10=0 $X=124660 $Y=48880 $D=28
M2714 VSS 3194 3205 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.37538e-14 as=2e-14 pd=4.70769e-07 ps=4e-07 nrd=1.09385 nrs=0.5 sa=6.8e-07 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=8.4e-15 panw7=1.56e-14 panw8=0 panw9=0 panw10=0 $X=124980 $Y=48880 $D=28
M2715 3206 543 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.79391e-13 pd=1.02e-06 ps=1.93015e-06 nrd=0.121951 nrs=0.266792 sa=4.49756e-07 sb=1.43244e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=125420 $Y=48390 $D=28
M2716 3194 3193 3206 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=7.69756e-07 sb=1.11244e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=125740 $Y=48390 $D=28
M2717 3207 3193 3194 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.24976e-06 sb=6.32439e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=126220 $Y=48390 $D=28
M2718 VSS 543 3207 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.47342e-13 as=8.2e-14 pd=2.16182e-06 ps=1.02e-06 nrd=0.367849 nrs=0.121951 sa=1.51122e-06 sb=3.12439e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=126540 $Y=48390 $D=28
M2719 3194 3196 3198 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.368e-13 pd=1.1e-06 ps=2.12e-06 nrd=0.243243 nrs=0.432432 sa=3.2e-07 sb=1.09189e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=127460 $Y=48710 $D=28
M2720 3198 3196 3194 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80119e-13 as=1.332e-13 pd=1.79489e-06 ps=1.1e-06 nrd=0.328925 nrs=0.243243 sa=8e-07 sb=6.33514e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=127940 $Y=48710 $D=28
M2721 3208 3195 3198 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=4.86809e-14 pd=4e-07 ps=4.85106e-07 nrd=0.5 nrs=1.21702 sa=1.32e-06 sb=1.08e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=128460 $Y=49050 $D=28
M2722 3209 543 3208 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.64e-06 sb=7.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=128780 $Y=49050 $D=28
M2723 VSS 3197 3209 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45167e-13 as=2e-14 pd=1.30833e-06 ps=4e-07 nrd=3.62917 nrs=0.5 sa=1.96e-06 sb=4.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=129100 $Y=49050 $D=28
M2724 VSS 3198 3197 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.87429e-14 as=9.84e-14 pd=4.65714e-07 ps=1.32e-06 nrd=1.21857 nrs=2.46 sa=3.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=130480 $Y=49110 $D=28
M2725 456 3198 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.24217e-13 pd=1.28e-06 ps=2.14229e-06 nrd=0.195652 nrs=0.264907 sa=3.97391e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=130880 $Y=48390 $D=28
M2726 VSS 3198 456 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8.77391e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=131360 $Y=48390 $D=28
M2727 VSS clk 3211 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.624e-13 as=1.792e-13 pd=1.28121e-06 ps=1.76e-06 nrd=0.517857 nrs=0.571429 sa=3.2e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=140410 $Y=41430 $D=28
M2728 3215 clk VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=1.392e-13 pd=1.68e-06 ps=1.09818e-06 nrd=0.75 nrs=0.604167 sa=8.8e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=140970 $Y=41510 $D=28
M2729 VSS 540 3212 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37856e-13 as=1.536e-13 pd=1.0432e-06 ps=1.6e-06 nrd=0.598333 nrs=0.666667 sa=3.2e-07 sb=1.10333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=142100 $Y=41630 $D=28
M2730 3216 3211 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.12528e-13 pd=2.6e-06 ps=1.60827e-06 nrd=0.588751 nrs=0.388108 sa=6.97297e-07 sb=4.35676e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=142660 $Y=41370 $D=28
M2731 3221 3215 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7e-14 as=2.88e-13 pd=9e-07 ps=2.54e-06 nrd=0.142857 nrs=0.587755 sa=3.27429e-07 sb=1.36e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=143840 $Y=41510 $D=28
M2732 3213 3212 3221 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=7e-14 pd=1.06e-06 ps=9e-07 nrd=0.257143 nrs=0.142857 sa=6.47429e-07 sb=1.04e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=144160 $Y=41510 $D=28
M2733 3223 3212 3213 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7e-14 as=1.26e-13 pd=9e-07 ps=1.06e-06 nrd=0.142857 nrs=0.257143 sa=1.12743e-06 sb=5.6e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=144640 $Y=41510 $D=28
M2734 VSS 3215 3223 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.32857e-13 as=7e-14 pd=2.35714e-06 ps=9e-07 nrd=0.475219 nrs=0.142857 sa=1.44743e-06 sb=2.4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=144960 $Y=41510 $D=28
M2735 3225 3216 3213 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=8.4e-15 panw7=1.56e-14 panw8=0 panw9=0 panw10=0 $X=145860 $Y=41680 $D=28
M2736 VSS 3214 3225 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.37538e-14 as=2e-14 pd=4.70769e-07 ps=4e-07 nrd=1.09385 nrs=0.5 sa=6.8e-07 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=8.4e-15 panw7=1.56e-14 panw8=0 panw9=0 panw10=0 $X=146180 $Y=41680 $D=28
M2737 3226 564 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.79391e-13 pd=1.02e-06 ps=1.93015e-06 nrd=0.121951 nrs=0.266792 sa=4.49756e-07 sb=1.43244e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=146620 $Y=41190 $D=28
M2738 3214 3213 3226 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=7.69756e-07 sb=1.11244e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=146940 $Y=41190 $D=28
M2739 3227 3213 3214 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.24976e-06 sb=6.32439e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=147420 $Y=41190 $D=28
M2740 VSS 564 3227 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.47342e-13 as=8.2e-14 pd=2.16182e-06 ps=1.02e-06 nrd=0.367849 nrs=0.121951 sa=1.51122e-06 sb=3.12439e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=147740 $Y=41190 $D=28
M2741 3214 3216 3218 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.368e-13 pd=1.1e-06 ps=2.12e-06 nrd=0.243243 nrs=0.432432 sa=3.2e-07 sb=1.09189e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=148660 $Y=41510 $D=28
M2742 3218 3216 3214 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80119e-13 as=1.332e-13 pd=1.79489e-06 ps=1.1e-06 nrd=0.328925 nrs=0.243243 sa=8e-07 sb=6.33514e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=149140 $Y=41510 $D=28
M2743 3228 3215 3218 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=4.86809e-14 pd=4e-07 ps=4.85106e-07 nrd=0.5 nrs=1.21702 sa=1.32e-06 sb=1.08e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=149660 $Y=41850 $D=28
M2744 3229 564 3228 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.64e-06 sb=7.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=149980 $Y=41850 $D=28
M2745 VSS 3217 3229 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45167e-13 as=2e-14 pd=1.30833e-06 ps=4e-07 nrd=3.62917 nrs=0.5 sa=1.96e-06 sb=4.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=150300 $Y=41850 $D=28
M2746 VSS 3218 3217 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.87429e-14 as=9.84e-14 pd=4.65714e-07 ps=1.32e-06 nrd=1.21857 nrs=2.46 sa=3.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=151680 $Y=41910 $D=28
M2747 568 3218 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.24217e-13 pd=1.28e-06 ps=2.14229e-06 nrd=0.195652 nrs=0.264907 sa=3.97391e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=152080 $Y=41190 $D=28
M2748 VSS 3218 568 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8.77391e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=152560 $Y=41190 $D=28
M2749 VSS clk 3231 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.624e-13 as=1.792e-13 pd=1.28121e-06 ps=1.76e-06 nrd=0.517857 nrs=0.571429 sa=3.2e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=146810 $Y=75610 $D=28
M2750 3235 clk VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=1.392e-13 pd=1.68e-06 ps=1.09818e-06 nrd=0.75 nrs=0.604167 sa=8.8e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=147370 $Y=75610 $D=28
M2751 VSS 856 3232 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37856e-13 as=1.536e-13 pd=1.0432e-06 ps=1.6e-06 nrd=0.598333 nrs=0.666667 sa=3.2e-07 sb=1.10333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=148500 $Y=75490 $D=28
M2752 3236 3231 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.12528e-13 pd=2.6e-06 ps=1.60827e-06 nrd=0.588751 nrs=0.388108 sa=6.97297e-07 sb=4.35676e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=149060 $Y=75490 $D=28
M2753 3241 3235 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7e-14 as=2.88e-13 pd=9e-07 ps=2.54e-06 nrd=0.142857 nrs=0.587755 sa=3.27429e-07 sb=1.36e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=150240 $Y=75390 $D=28
M2754 3233 3232 3241 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=7e-14 pd=1.06e-06 ps=9e-07 nrd=0.257143 nrs=0.142857 sa=6.47429e-07 sb=1.04e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=150560 $Y=75390 $D=28
M2755 3243 3232 3233 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7e-14 as=1.26e-13 pd=9e-07 ps=1.06e-06 nrd=0.142857 nrs=0.257143 sa=1.12743e-06 sb=5.6e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=151040 $Y=75390 $D=28
M2756 VSS 3235 3243 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.32857e-13 as=7e-14 pd=2.35714e-06 ps=9e-07 nrd=0.475219 nrs=0.142857 sa=1.44743e-06 sb=2.4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=151360 $Y=75390 $D=28
M2757 3245 3236 3233 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=8.4e-15 panw7=1.56e-14 panw8=0 panw9=0 panw10=0 $X=152260 $Y=75720 $D=28
M2758 VSS 3234 3245 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.37538e-14 as=2e-14 pd=4.70769e-07 ps=4e-07 nrd=1.09385 nrs=0.5 sa=6.8e-07 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=8.4e-15 panw7=1.56e-14 panw8=0 panw9=0 panw10=0 $X=152580 $Y=75720 $D=28
M2759 3246 610 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.79391e-13 pd=1.02e-06 ps=1.93015e-06 nrd=0.121951 nrs=0.266792 sa=4.49756e-07 sb=1.43244e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=153020 $Y=75590 $D=28
M2760 3234 3233 3246 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=7.69756e-07 sb=1.11244e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=153340 $Y=75590 $D=28
M2761 3247 3233 3234 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.24976e-06 sb=6.32439e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=153820 $Y=75590 $D=28
M2762 VSS 610 3247 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.47342e-13 as=8.2e-14 pd=2.16182e-06 ps=1.02e-06 nrd=0.367849 nrs=0.121951 sa=1.51122e-06 sb=3.12439e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=154140 $Y=75590 $D=28
M2763 3234 3236 3238 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.368e-13 pd=1.1e-06 ps=2.12e-06 nrd=0.243243 nrs=0.432432 sa=3.2e-07 sb=1.09189e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=155060 $Y=75350 $D=28
M2764 3238 3236 3234 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80119e-13 as=1.332e-13 pd=1.79489e-06 ps=1.1e-06 nrd=0.328925 nrs=0.243243 sa=8e-07 sb=6.33514e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=155540 $Y=75350 $D=28
M2765 3248 3235 3238 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=4.86809e-14 pd=4e-07 ps=4.85106e-07 nrd=0.5 nrs=1.21702 sa=1.32e-06 sb=1.08e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=156060 $Y=75550 $D=28
M2766 3249 610 3248 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.64e-06 sb=7.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=156380 $Y=75550 $D=28
M2767 VSS 3237 3249 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45167e-13 as=2e-14 pd=1.30833e-06 ps=4e-07 nrd=3.62917 nrs=0.5 sa=1.96e-06 sb=4.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=156700 $Y=75550 $D=28
M2768 VSS 3238 3237 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.87429e-14 as=9.84e-14 pd=4.65714e-07 ps=1.32e-06 nrd=1.21857 nrs=2.46 sa=3.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=158080 $Y=75490 $D=28
M2769 609 3238 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.24217e-13 pd=1.28e-06 ps=2.14229e-06 nrd=0.195652 nrs=0.264907 sa=3.97391e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=158480 $Y=75490 $D=28
M2770 VSS 3238 609 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8.77391e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=158960 $Y=75490 $D=28
M2771 VSS clk 3251 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.624e-13 as=1.792e-13 pd=1.28121e-06 ps=1.76e-06 nrd=0.517857 nrs=0.571429 sa=3.2e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=164810 $Y=54010 $D=28
M2772 3255 clk VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=1.392e-13 pd=1.68e-06 ps=1.09818e-06 nrd=0.75 nrs=0.604167 sa=8.8e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=165370 $Y=54010 $D=28
M2773 VSS 664 3252 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37856e-13 as=1.536e-13 pd=1.0432e-06 ps=1.6e-06 nrd=0.598333 nrs=0.666667 sa=3.2e-07 sb=1.10333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=166500 $Y=53890 $D=28
M2774 3256 3251 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.12528e-13 pd=2.6e-06 ps=1.60827e-06 nrd=0.588751 nrs=0.388108 sa=6.97297e-07 sb=4.35676e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=167060 $Y=53890 $D=28
M2775 3261 3255 VSS VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7e-14 as=2.88e-13 pd=9e-07 ps=2.54e-06 nrd=0.142857 nrs=0.587755 sa=3.27429e-07 sb=1.36e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=168240 $Y=53790 $D=28
M2776 3253 3252 3261 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=7e-14 pd=1.06e-06 ps=9e-07 nrd=0.257143 nrs=0.142857 sa=6.47429e-07 sb=1.04e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=168560 $Y=53790 $D=28
M2777 3263 3252 3253 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7e-14 as=1.26e-13 pd=9e-07 ps=1.06e-06 nrd=0.142857 nrs=0.257143 sa=1.12743e-06 sb=5.6e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=169040 $Y=53790 $D=28
M2778 VSS 3255 3263 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.32857e-13 as=7e-14 pd=2.35714e-06 ps=9e-07 nrd=0.475219 nrs=0.142857 sa=1.44743e-06 sb=2.4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-15 panw10=0 $X=169360 $Y=53790 $D=28
M2779 3265 3256 3253 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=8.4e-15 panw7=1.56e-14 panw8=0 panw9=0 panw10=0 $X=170260 $Y=54120 $D=28
M2780 VSS 3254 3265 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.37538e-14 as=2e-14 pd=4.70769e-07 ps=4e-07 nrd=1.09385 nrs=0.5 sa=6.8e-07 sb=1.86e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=8.4e-15 panw7=1.56e-14 panw8=0 panw9=0 panw10=0 $X=170580 $Y=54120 $D=28
M2781 3266 697 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.79391e-13 pd=1.02e-06 ps=1.93015e-06 nrd=0.121951 nrs=0.266792 sa=4.49756e-07 sb=1.43244e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=171020 $Y=53990 $D=28
M2782 3254 3253 3266 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=7.69756e-07 sb=1.11244e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=171340 $Y=53990 $D=28
M2783 3267 3253 3254 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.24976e-06 sb=6.32439e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=171820 $Y=53990 $D=28
M2784 VSS 697 3267 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.47342e-13 as=8.2e-14 pd=2.16182e-06 ps=1.02e-06 nrd=0.367849 nrs=0.121951 sa=1.51122e-06 sb=3.12439e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=172140 $Y=53990 $D=28
M2785 3254 3256 3258 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.368e-13 pd=1.1e-06 ps=2.12e-06 nrd=0.243243 nrs=0.432432 sa=3.2e-07 sb=1.09189e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=173060 $Y=53750 $D=28
M2786 3258 3256 3254 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80119e-13 as=1.332e-13 pd=1.79489e-06 ps=1.1e-06 nrd=0.328925 nrs=0.243243 sa=8e-07 sb=6.33514e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=173540 $Y=53750 $D=28
M2787 3268 3255 3258 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=4.86809e-14 pd=4e-07 ps=4.85106e-07 nrd=0.5 nrs=1.21702 sa=1.32e-06 sb=1.08e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=174060 $Y=53950 $D=28
M2788 3269 697 3268 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=1.64e-06 sb=7.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=174380 $Y=53950 $D=28
M2789 VSS 3257 3269 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45167e-13 as=2e-14 pd=1.30833e-06 ps=4e-07 nrd=3.62917 nrs=0.5 sa=1.96e-06 sb=4.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=174700 $Y=53950 $D=28
M2790 VSS 3258 3257 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.87429e-14 as=9.84e-14 pd=4.65714e-07 ps=1.32e-06 nrd=1.21857 nrs=2.46 sa=3.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=176080 $Y=53890 $D=28
M2791 597 3258 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.24217e-13 pd=1.28e-06 ps=2.14229e-06 nrd=0.195652 nrs=0.264907 sa=3.97391e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=176480 $Y=53890 $D=28
M2792 VSS 3258 597 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8.77391e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=176960 $Y=53890 $D=28
M2793 VSS data_in[5] 3271 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=8860 $Y=53890 $D=28
M2794 157 3271 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=9440 $Y=53890 $D=28
M2795 VSS 797 3272 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=10460 $Y=53890 $D=28
M2796 183 3272 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=11040 $Y=53890 $D=28
M2797 VSS 318 3273 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=86460 $Y=25090 $D=28
M2798 300 3273 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=87040 $Y=25090 $D=28
M2799 VSS 306 3274 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=88060 $Y=25090 $D=28
M2800 345 3274 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=88640 $Y=25090 $D=28
M2801 VSS 377 3275 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=92860 $Y=20310 $D=28
M2802 318 3275 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=93440 $Y=20030 $D=28
M2803 VSS 345 3276 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=94460 $Y=20310 $D=28
M2804 368 3276 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=95040 $Y=20030 $D=28
M2805 VSS 329 3277 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=98460 $Y=27510 $D=28
M2806 407 3277 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=99040 $Y=27230 $D=28
M2807 VSS 377 3278 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=100060 $Y=27510 $D=28
M2808 409 3278 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=100640 $Y=27230 $D=28
M2809 VSS 377 3279 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=102860 $Y=20310 $D=28
M2810 399 3279 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=103440 $Y=20030 $D=28
M2811 VSS 368 3280 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=104460 $Y=20310 $D=28
M2812 396 3280 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=105040 $Y=20030 $D=28
M2813 VSS 390 3281 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=106060 $Y=20310 $D=28
M2814 data_out[0] 3281 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=106640 $Y=20030 $D=28
M2815 VSS 399 3282 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=107660 $Y=20310 $D=28
M2816 408 3282 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=108240 $Y=20030 $D=28
M2817 VSS 543 3283 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=141660 $Y=49110 $D=28
M2818 544 3283 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=142240 $Y=48830 $D=28
M2819 VSS 544 3284 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=143260 $Y=49110 $D=28
M2820 697 3284 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=143840 $Y=48830 $D=28
M2821 VSS 611 3285 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=153260 $Y=20310 $D=28
M2822 682 3285 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=153840 $Y=20030 $D=28
M2823 VSS 570 3286 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.83529e-14 as=9.44e-14 pd=5.52941e-07 ps=1.28e-06 nrd=1.45882 nrs=2.36 sa=3.6e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=154860 $Y=20310 $D=28
M2824 620 3286 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=1.40047e-13 pd=1.6e-06 ps=1.32706e-06 nrd=0.666667 nrs=0.607843 sa=6.13333e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=155440 $Y=20030 $D=28
M2825 3296 3289 3290 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=11660 $Y=10710 $D=28
M2826 3298 97 3296 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=11980 $Y=10710 $D=28
M2827 VSS 76 3298 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=12300 $Y=10710 $D=28
M2828 VSS clk 3289 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=13280 $Y=10860 $D=28
M2829 3292 3289 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=13790 $Y=10860 $D=28
M2830 3300 3292 3290 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=14810 $Y=10790 $D=28
M2831 3301 3291 3300 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=15130 $Y=10790 $D=28
M2832 VSS 76 3301 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=15450 $Y=10790 $D=28
M2833 3291 3290 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=15910 $Y=10930 $D=28
M2834 3293 3292 3291 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=16470 $Y=10930 $D=28
M2835 3303 3289 3293 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=17030 $Y=10690 $D=28
M2836 VSS 3295 3303 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=17350 $Y=10690 $D=28
M2837 3304 76 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=17790 $Y=10690 $D=28
M2838 3295 3293 3304 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=18110 $Y=10690 $D=28
M2839 3294 3295 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=18430 $Y=11410 $D=28
M2840 VSS 3294 3287 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=19330 $Y=10690 $D=28
M2841 weight_out[0] 3295 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=19830 $Y=10690 $D=28
M2842 3312 3305 3306 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=20860 $Y=10710 $D=28
M2843 3314 79 3312 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=21180 $Y=10710 $D=28
M2844 VSS 76 3314 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=21500 $Y=10710 $D=28
M2845 VSS clk 3305 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=22480 $Y=10860 $D=28
M2846 3308 3305 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=22990 $Y=10860 $D=28
M2847 3316 3308 3306 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=24010 $Y=10790 $D=28
M2848 3317 3307 3316 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=24330 $Y=10790 $D=28
M2849 VSS 76 3317 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=24650 $Y=10790 $D=28
M2850 3307 3306 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=25110 $Y=10930 $D=28
M2851 3309 3308 3307 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=25670 $Y=10930 $D=28
M2852 3319 3305 3309 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=26230 $Y=10690 $D=28
M2853 VSS 3311 3319 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=26550 $Y=10690 $D=28
M2854 3320 76 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=26990 $Y=10690 $D=28
M2855 3311 3309 3320 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=27310 $Y=10690 $D=28
M2856 3310 3311 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=27630 $Y=11410 $D=28
M2857 VSS 3310 3288 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=28530 $Y=10690 $D=28
M2858 weight_out[2] 3311 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=29030 $Y=10690 $D=28
M2859 3330 3323 3324 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=30060 $Y=10710 $D=28
M2860 3332 113 3330 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=30380 $Y=10710 $D=28
M2861 VSS 128 3332 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=30700 $Y=10710 $D=28
M2862 VSS clk 3323 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=31680 $Y=10860 $D=28
M2863 3326 3323 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=32190 $Y=10860 $D=28
M2864 3334 3326 3324 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=33210 $Y=10790 $D=28
M2865 3335 3325 3334 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=33530 $Y=10790 $D=28
M2866 VSS 128 3335 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=33850 $Y=10790 $D=28
M2867 3325 3324 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=34310 $Y=10930 $D=28
M2868 3327 3326 3325 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=34870 $Y=10930 $D=28
M2869 3337 3323 3327 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=35430 $Y=10690 $D=28
M2870 VSS 3329 3337 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=35750 $Y=10690 $D=28
M2871 3338 128 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=36190 $Y=10690 $D=28
M2872 3329 3327 3338 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=36510 $Y=10690 $D=28
M2873 3328 3329 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=36830 $Y=11410 $D=28
M2874 VSS 3328 3321 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=37730 $Y=10690 $D=28
M2875 weight_out[1] 3329 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=38230 $Y=10690 $D=28
M2876 3346 3339 3340 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=39260 $Y=10710 $D=28
M2877 3348 195 3346 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=39580 $Y=10710 $D=28
M2878 VSS 202 3348 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=39900 $Y=10710 $D=28
M2879 VSS clk 3339 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=40880 $Y=10860 $D=28
M2880 3342 3339 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=41390 $Y=10860 $D=28
M2881 3350 3342 3340 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=42410 $Y=10790 $D=28
M2882 3351 3341 3350 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=42730 $Y=10790 $D=28
M2883 VSS 202 3351 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=43050 $Y=10790 $D=28
M2884 3341 3340 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=43510 $Y=10930 $D=28
M2885 3343 3342 3341 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=44070 $Y=10930 $D=28
M2886 3353 3339 3343 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=44630 $Y=10690 $D=28
M2887 VSS 3345 3353 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=44950 $Y=10690 $D=28
M2888 3354 202 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=45390 $Y=10690 $D=28
M2889 3345 3343 3354 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=45710 $Y=10690 $D=28
M2890 3344 3345 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=46030 $Y=11410 $D=28
M2891 VSS 3344 3322 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=46930 $Y=10690 $D=28
M2892 weight_out[6] 3345 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=47430 $Y=10690 $D=28
M2893 3364 3357 3358 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=36060 $Y=13090 $D=28
M2894 3366 135 3364 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=36380 $Y=13090 $D=28
M2895 VSS 128 3366 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=36700 $Y=13090 $D=28
M2896 VSS clk 3357 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=37680 $Y=12840 $D=28
M2897 3360 3357 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=38190 $Y=12940 $D=28
M2898 3368 3360 3358 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=39210 $Y=13010 $D=28
M2899 3369 3359 3368 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=39530 $Y=13010 $D=28
M2900 VSS 128 3369 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=39850 $Y=13010 $D=28
M2901 3359 3358 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=40310 $Y=12870 $D=28
M2902 3361 3360 3359 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=40870 $Y=12870 $D=28
M2903 3371 3357 3361 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=41430 $Y=13110 $D=28
M2904 VSS 3363 3371 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=41750 $Y=13110 $D=28
M2905 3372 128 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=42190 $Y=13090 $D=28
M2906 3363 3361 3372 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=42510 $Y=13090 $D=28
M2907 3362 3363 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=42830 $Y=12390 $D=28
M2908 VSS 3362 3355 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=43730 $Y=13070 $D=28
M2909 weight_out[4] 3363 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=44230 $Y=13070 $D=28
M2910 3380 3373 3374 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=45260 $Y=13090 $D=28
M2911 3382 170 3380 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=45580 $Y=13090 $D=28
M2912 VSS 128 3382 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=45900 $Y=13090 $D=28
M2913 VSS clk 3373 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=46880 $Y=12840 $D=28
M2914 3376 3373 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=47390 $Y=12940 $D=28
M2915 3384 3376 3374 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=48410 $Y=13010 $D=28
M2916 3385 3375 3384 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=48730 $Y=13010 $D=28
M2917 VSS 128 3385 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=49050 $Y=13010 $D=28
M2918 3375 3374 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=49510 $Y=12870 $D=28
M2919 3377 3376 3375 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=50070 $Y=12870 $D=28
M2920 3387 3373 3377 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=50630 $Y=13110 $D=28
M2921 VSS 3379 3387 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=50950 $Y=13110 $D=28
M2922 3388 128 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=51390 $Y=13090 $D=28
M2923 3379 3377 3388 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=51710 $Y=13090 $D=28
M2924 3378 3379 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=52030 $Y=12390 $D=28
M2925 VSS 3378 3356 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=52930 $Y=13070 $D=28
M2926 weight_out[5] 3379 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=53430 $Y=13070 $D=28
M2927 3398 3391 3392 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=50460 $Y=10710 $D=28
M2928 3400 240 3398 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=50780 $Y=10710 $D=28
M2929 VSS 202 3400 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=51100 $Y=10710 $D=28
M2930 VSS clk 3391 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=52080 $Y=10860 $D=28
M2931 3394 3391 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=52590 $Y=10860 $D=28
M2932 3402 3394 3392 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=53610 $Y=10790 $D=28
M2933 3403 3393 3402 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=53930 $Y=10790 $D=28
M2934 VSS 202 3403 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=54250 $Y=10790 $D=28
M2935 3393 3392 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=54710 $Y=10930 $D=28
M2936 3395 3394 3393 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=55270 $Y=10930 $D=28
M2937 3405 3391 3395 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=55830 $Y=10690 $D=28
M2938 VSS 3397 3405 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=56150 $Y=10690 $D=28
M2939 3406 202 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=56590 $Y=10690 $D=28
M2940 3397 3395 3406 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=56910 $Y=10690 $D=28
M2941 3396 3397 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=57230 $Y=11410 $D=28
M2942 VSS 3396 3389 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=58130 $Y=10690 $D=28
M2943 weight_out[7] 3397 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=58630 $Y=10690 $D=28
M2944 3414 3407 3408 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=59660 $Y=10710 $D=28
M2945 3416 310 3414 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=59980 $Y=10710 $D=28
M2946 VSS 252 3416 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=60300 $Y=10710 $D=28
M2947 VSS clk 3407 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=61280 $Y=10860 $D=28
M2948 3410 3407 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=61790 $Y=10860 $D=28
M2949 3418 3410 3408 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=62810 $Y=10790 $D=28
M2950 3419 3409 3418 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=63130 $Y=10790 $D=28
M2951 VSS 252 3419 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=63450 $Y=10790 $D=28
M2952 3409 3408 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=63910 $Y=10930 $D=28
M2953 3411 3410 3409 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=64470 $Y=10930 $D=28
M2954 3421 3407 3411 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=65030 $Y=10690 $D=28
M2955 VSS 3413 3421 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=65350 $Y=10690 $D=28
M2956 3422 252 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=65790 $Y=10690 $D=28
M2957 3413 3411 3422 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=66110 $Y=10690 $D=28
M2958 3412 3413 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=66430 $Y=11410 $D=28
M2959 VSS 3412 3390 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=67330 $Y=10690 $D=28
M2960 fire_out 3413 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=67830 $Y=10690 $D=28
M2961 3432 3425 3426 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=68860 $Y=10710 $D=28
M2962 3434 251 3432 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=69180 $Y=10710 $D=28
M2963 VSS 252 3434 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=69500 $Y=10710 $D=28
M2964 VSS clk 3425 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=70480 $Y=10860 $D=28
M2965 3428 3425 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=70990 $Y=10860 $D=28
M2966 3436 3428 3426 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=72010 $Y=10790 $D=28
M2967 3437 3427 3436 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=72330 $Y=10790 $D=28
M2968 VSS 252 3437 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=72650 $Y=10790 $D=28
M2969 3427 3426 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=73110 $Y=10930 $D=28
M2970 3429 3428 3427 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=73670 $Y=10930 $D=28
M2971 3439 3425 3429 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=74230 $Y=10690 $D=28
M2972 VSS 3431 3439 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=74550 $Y=10690 $D=28
M2973 3440 252 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=74990 $Y=10690 $D=28
M2974 3431 3429 3440 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=75310 $Y=10690 $D=28
M2975 3430 3431 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=75630 $Y=11410 $D=28
M2976 VSS 3430 3423 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=76530 $Y=10690 $D=28
M2977 result[1] 3431 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=77030 $Y=10690 $D=28
M2978 3448 3441 3442 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=78060 $Y=10710 $D=28
M2979 3450 828 3448 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=78380 $Y=10710 $D=28
M2980 VSS 299 3450 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=78700 $Y=10710 $D=28
M2981 VSS clk 3441 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=79680 $Y=10860 $D=28
M2982 3444 3441 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=80190 $Y=10860 $D=28
M2983 3452 3444 3442 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=81210 $Y=10790 $D=28
M2984 3453 3443 3452 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=81530 $Y=10790 $D=28
M2985 VSS 299 3453 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=81850 $Y=10790 $D=28
M2986 3443 3442 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=82310 $Y=10930 $D=28
M2987 3445 3444 3443 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=82870 $Y=10930 $D=28
M2988 3455 3441 3445 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=83430 $Y=10690 $D=28
M2989 VSS 3447 3455 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=83750 $Y=10690 $D=28
M2990 3456 299 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=84190 $Y=10690 $D=28
M2991 3447 3445 3456 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=84510 $Y=10690 $D=28
M2992 3446 3447 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=84830 $Y=11410 $D=28
M2993 VSS 3446 3424 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=85730 $Y=10690 $D=28
M2994 result[2] 3447 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=86230 $Y=10690 $D=28
M2995 3466 3459 3460 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=80060 $Y=27490 $D=28
M2996 3468 305 3466 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=80380 $Y=27490 $D=28
M2997 VSS 303 3468 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=80700 $Y=27490 $D=28
M2998 VSS clk 3459 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=81680 $Y=27240 $D=28
M2999 3462 3459 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=82190 $Y=27340 $D=28
M3000 3470 3462 3460 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=83210 $Y=27410 $D=28
M3001 3471 3461 3470 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=83530 $Y=27410 $D=28
M3002 VSS 303 3471 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=83850 $Y=27410 $D=28
M3003 3461 3460 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=84310 $Y=27270 $D=28
M3004 3463 3462 3461 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=84870 $Y=27270 $D=28
M3005 3473 3459 3463 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=85430 $Y=27510 $D=28
M3006 VSS 3465 3473 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=85750 $Y=27510 $D=28
M3007 3474 303 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=86190 $Y=27490 $D=28
M3008 3465 3463 3474 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=86510 $Y=27490 $D=28
M3009 3464 3465 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=86830 $Y=26790 $D=28
M3010 VSS 3464 3457 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=87730 $Y=27470 $D=28
M3011 result[5] 3465 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=88230 $Y=27470 $D=28
M3012 3482 3475 3476 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=89260 $Y=27490 $D=28
M3013 3484 217 3482 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=89580 $Y=27490 $D=28
M3014 VSS 329 3484 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=89900 $Y=27490 $D=28
M3015 VSS clk 3475 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=90880 $Y=27240 $D=28
M3016 3478 3475 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=91390 $Y=27340 $D=28
M3017 3486 3478 3476 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=92410 $Y=27410 $D=28
M3018 3487 3477 3486 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=92730 $Y=27410 $D=28
M3019 VSS 329 3487 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=93050 $Y=27410 $D=28
M3020 3477 3476 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=93510 $Y=27270 $D=28
M3021 3479 3478 3477 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=94070 $Y=27270 $D=28
M3022 3489 3475 3479 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=94630 $Y=27510 $D=28
M3023 VSS 3481 3489 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=94950 $Y=27510 $D=28
M3024 3490 329 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=95390 $Y=27490 $D=28
M3025 3481 3479 3490 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=95710 $Y=27490 $D=28
M3026 3480 3481 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=96030 $Y=26790 $D=28
M3027 VSS 3480 3458 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96930 $Y=27470 $D=28
M3028 390 3481 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=97430 $Y=27470 $D=28
M3029 3500 3493 3494 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=87260 $Y=10710 $D=28
M3030 3502 333 3500 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=87580 $Y=10710 $D=28
M3031 VSS 356 3502 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=87900 $Y=10710 $D=28
M3032 VSS clk 3493 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=88880 $Y=10860 $D=28
M3033 3496 3493 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=89390 $Y=10860 $D=28
M3034 3504 3496 3494 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=90410 $Y=10790 $D=28
M3035 3505 3495 3504 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=90730 $Y=10790 $D=28
M3036 VSS 356 3505 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=91050 $Y=10790 $D=28
M3037 3495 3494 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=91510 $Y=10930 $D=28
M3038 3497 3496 3495 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=92070 $Y=10930 $D=28
M3039 3507 3493 3497 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=92630 $Y=10690 $D=28
M3040 VSS 3499 3507 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=92950 $Y=10690 $D=28
M3041 3508 356 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=93390 $Y=10690 $D=28
M3042 3499 3497 3508 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=93710 $Y=10690 $D=28
M3043 3498 3499 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=94030 $Y=11410 $D=28
M3044 VSS 3498 3491 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=94930 $Y=10690 $D=28
M3045 result[3] 3499 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=95430 $Y=10690 $D=28
M3046 3516 3509 3510 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96460 $Y=10710 $D=28
M3047 3518 364 3516 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96780 $Y=10710 $D=28
M3048 VSS 356 3518 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=97100 $Y=10710 $D=28
M3049 VSS clk 3509 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=98080 $Y=10860 $D=28
M3050 3512 3509 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=98590 $Y=10860 $D=28
M3051 3520 3512 3510 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=99610 $Y=10790 $D=28
M3052 3521 3511 3520 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=99930 $Y=10790 $D=28
M3053 VSS 356 3521 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=100250 $Y=10790 $D=28
M3054 3511 3510 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=100710 $Y=10930 $D=28
M3055 3513 3512 3511 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=101270 $Y=10930 $D=28
M3056 3523 3509 3513 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=101830 $Y=10690 $D=28
M3057 VSS 3515 3523 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=102150 $Y=10690 $D=28
M3058 3524 356 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=102590 $Y=10690 $D=28
M3059 3515 3513 3524 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=102910 $Y=10690 $D=28
M3060 3514 3515 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=103230 $Y=11410 $D=28
M3061 VSS 3514 3492 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=104130 $Y=10690 $D=28
M3062 result[10] 3515 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=104630 $Y=10690 $D=28
M3063 3534 3527 3528 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=89660 $Y=25110 $D=28
M3064 3536 332 3534 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=89980 $Y=25110 $D=28
M3065 VSS 329 3536 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=90300 $Y=25110 $D=28
M3066 VSS clk 3527 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=91280 $Y=25260 $D=28
M3067 3530 3527 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=91790 $Y=25260 $D=28
M3068 3538 3530 3528 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=92810 $Y=25190 $D=28
M3069 3539 3529 3538 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=93130 $Y=25190 $D=28
M3070 VSS 329 3539 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=93450 $Y=25190 $D=28
M3071 3529 3528 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=93910 $Y=25330 $D=28
M3072 3531 3530 3529 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=94470 $Y=25330 $D=28
M3073 3541 3527 3531 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=95030 $Y=25090 $D=28
M3074 VSS 3533 3541 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=95350 $Y=25090 $D=28
M3075 3542 329 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=95790 $Y=25090 $D=28
M3076 3533 3531 3542 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96110 $Y=25090 $D=28
M3077 3532 3533 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=96430 $Y=25810 $D=28
M3078 VSS 3532 3525 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=97330 $Y=25090 $D=28
M3079 result[7] 3533 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=97830 $Y=25090 $D=28
M3080 3550 3543 3544 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=98860 $Y=25110 $D=28
M3081 3552 832 3550 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=99180 $Y=25110 $D=28
M3082 VSS 407 3552 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=99500 $Y=25110 $D=28
M3083 VSS clk 3543 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=100480 $Y=25260 $D=28
M3084 3546 3543 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=100990 $Y=25260 $D=28
M3085 3554 3546 3544 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=102010 $Y=25190 $D=28
M3086 3555 3545 3554 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=102330 $Y=25190 $D=28
M3087 VSS 407 3555 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=102650 $Y=25190 $D=28
M3088 3545 3544 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=103110 $Y=25330 $D=28
M3089 3547 3546 3545 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=103670 $Y=25330 $D=28
M3090 3557 3543 3547 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=104230 $Y=25090 $D=28
M3091 VSS 3549 3557 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=104550 $Y=25090 $D=28
M3092 3558 407 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=104990 $Y=25090 $D=28
M3093 3549 3547 3558 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=105310 $Y=25090 $D=28
M3094 3548 3549 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=105630 $Y=25810 $D=28
M3095 VSS 3548 3526 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=106530 $Y=25090 $D=28
M3096 result[8] 3549 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=107030 $Y=25090 $D=28
M3097 3568 3561 3562 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=105260 $Y=13090 $D=28
M3098 3570 388 3568 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=105580 $Y=13090 $D=28
M3099 VSS 371 3570 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=105900 $Y=13090 $D=28
M3100 VSS clk 3561 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=106880 $Y=12840 $D=28
M3101 3564 3561 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=107390 $Y=12940 $D=28
M3102 3572 3564 3562 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=108410 $Y=13010 $D=28
M3103 3573 3563 3572 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=108730 $Y=13010 $D=28
M3104 VSS 371 3573 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=109050 $Y=13010 $D=28
M3105 3563 3562 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=109510 $Y=12870 $D=28
M3106 3565 3564 3563 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=110070 $Y=12870 $D=28
M3107 3575 3561 3565 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=110630 $Y=13110 $D=28
M3108 VSS 3567 3575 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=110950 $Y=13110 $D=28
M3109 3576 371 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=111390 $Y=13090 $D=28
M3110 3567 3565 3576 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=111710 $Y=13090 $D=28
M3111 3566 3567 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=112030 $Y=12390 $D=28
M3112 VSS 3566 3559 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=112930 $Y=13070 $D=28
M3113 result[12] 3567 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=113430 $Y=13070 $D=28
M3114 3584 3577 3578 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=114460 $Y=13090 $D=28
M3115 3586 424 3584 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=114780 $Y=13090 $D=28
M3116 VSS 428 3586 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=115100 $Y=13090 $D=28
M3117 VSS clk 3577 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=116080 $Y=12840 $D=28
M3118 3580 3577 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=116590 $Y=12940 $D=28
M3119 3588 3580 3578 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=117610 $Y=13010 $D=28
M3120 3589 3579 3588 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=117930 $Y=13010 $D=28
M3121 VSS 428 3589 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=118250 $Y=13010 $D=28
M3122 3579 3578 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=118710 $Y=12870 $D=28
M3123 3581 3580 3579 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=119270 $Y=12870 $D=28
M3124 3591 3577 3581 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=119830 $Y=13110 $D=28
M3125 VSS 3583 3591 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=120150 $Y=13110 $D=28
M3126 3592 428 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=120590 $Y=13090 $D=28
M3127 3583 3581 3592 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=120910 $Y=13090 $D=28
M3128 3582 3583 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=121230 $Y=12390 $D=28
M3129 VSS 3582 3560 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=122130 $Y=13070 $D=28
M3130 result[15] 3583 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=122630 $Y=13070 $D=28
M3131 3602 3595 3596 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=119260 $Y=10710 $D=28
M3132 3604 449 3602 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=119580 $Y=10710 $D=28
M3133 VSS 479 3604 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=119900 $Y=10710 $D=28
M3134 VSS clk 3595 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=120880 $Y=10860 $D=28
M3135 3598 3595 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=121390 $Y=10860 $D=28
M3136 3606 3598 3596 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=122410 $Y=10790 $D=28
M3137 3607 3597 3606 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=122730 $Y=10790 $D=28
M3138 VSS 479 3607 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=123050 $Y=10790 $D=28
M3139 3597 3596 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=123510 $Y=10930 $D=28
M3140 3599 3598 3597 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=124070 $Y=10930 $D=28
M3141 3609 3595 3599 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=124630 $Y=10690 $D=28
M3142 VSS 3601 3609 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=124950 $Y=10690 $D=28
M3143 3610 479 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=125390 $Y=10690 $D=28
M3144 3601 3599 3610 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=125710 $Y=10690 $D=28
M3145 3600 3601 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=126030 $Y=11410 $D=28
M3146 VSS 3600 3593 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=126930 $Y=10690 $D=28
M3147 result[16] 3601 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=127430 $Y=10690 $D=28
M3148 3618 3611 3612 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=128460 $Y=10710 $D=28
M3149 3620 513 3618 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=128780 $Y=10710 $D=28
M3150 VSS 479 3620 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=129100 $Y=10710 $D=28
M3151 VSS clk 3611 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=130080 $Y=10860 $D=28
M3152 3614 3611 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=130590 $Y=10860 $D=28
M3153 3622 3614 3612 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=131610 $Y=10790 $D=28
M3154 3623 3613 3622 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=131930 $Y=10790 $D=28
M3155 VSS 479 3623 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=132250 $Y=10790 $D=28
M3156 3613 3612 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=132710 $Y=10930 $D=28
M3157 3615 3614 3613 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=133270 $Y=10930 $D=28
M3158 3625 3611 3615 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=133830 $Y=10690 $D=28
M3159 VSS 3617 3625 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=134150 $Y=10690 $D=28
M3160 3626 479 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=134590 $Y=10690 $D=28
M3161 3617 3615 3626 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=134910 $Y=10690 $D=28
M3162 3616 3617 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=135230 $Y=11410 $D=28
M3163 VSS 3616 3594 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=136130 $Y=10690 $D=28
M3164 result[17] 3617 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=136630 $Y=10690 $D=28
M3165 3636 3629 3630 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=137660 $Y=10710 $D=28
M3166 3638 541 3636 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=137980 $Y=10710 $D=28
M3167 VSS 584 3638 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=138300 $Y=10710 $D=28
M3168 VSS clk 3629 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=139280 $Y=10860 $D=28
M3169 3632 3629 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=139790 $Y=10860 $D=28
M3170 3640 3632 3630 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=140810 $Y=10790 $D=28
M3171 3641 3631 3640 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=141130 $Y=10790 $D=28
M3172 VSS 584 3641 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=141450 $Y=10790 $D=28
M3173 3631 3630 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=141910 $Y=10930 $D=28
M3174 3633 3632 3631 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=142470 $Y=10930 $D=28
M3175 3643 3629 3633 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=143030 $Y=10690 $D=28
M3176 VSS 3635 3643 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=143350 $Y=10690 $D=28
M3177 3644 584 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=143790 $Y=10690 $D=28
M3178 3635 3633 3644 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=144110 $Y=10690 $D=28
M3179 3634 3635 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=144430 $Y=11410 $D=28
M3180 VSS 3634 3627 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=145330 $Y=10690 $D=28
M3181 result[18] 3635 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=145830 $Y=10690 $D=28
M3182 3652 3645 3646 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=146860 $Y=10710 $D=28
M3183 3654 604 3652 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=147180 $Y=10710 $D=28
M3184 VSS 584 3654 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=147500 $Y=10710 $D=28
M3185 VSS clk 3645 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=148480 $Y=10860 $D=28
M3186 3648 3645 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=148990 $Y=10860 $D=28
M3187 3656 3648 3646 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=150010 $Y=10790 $D=28
M3188 3657 3647 3656 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=150330 $Y=10790 $D=28
M3189 VSS 584 3657 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=150650 $Y=10790 $D=28
M3190 3647 3646 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=151110 $Y=10930 $D=28
M3191 3649 3648 3647 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=151670 $Y=10930 $D=28
M3192 3659 3645 3649 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=152230 $Y=10690 $D=28
M3193 VSS 3651 3659 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=152550 $Y=10690 $D=28
M3194 3660 584 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=152990 $Y=10690 $D=28
M3195 3651 3649 3660 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=153310 $Y=10690 $D=28
M3196 3650 3651 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=153630 $Y=11410 $D=28
M3197 VSS 3650 3628 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=154530 $Y=10690 $D=28
M3198 result[21] 3651 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=155030 $Y=10690 $D=28
M3199 3670 3663 3664 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=140860 $Y=13090 $D=28
M3200 3672 579 3670 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=141180 $Y=13090 $D=28
M3201 VSS 584 3672 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=141500 $Y=13090 $D=28
M3202 VSS clk 3663 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=142480 $Y=12840 $D=28
M3203 3666 3663 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=142990 $Y=12940 $D=28
M3204 3674 3666 3664 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=144010 $Y=13010 $D=28
M3205 3675 3665 3674 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=144330 $Y=13010 $D=28
M3206 VSS 584 3675 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=144650 $Y=13010 $D=28
M3207 3665 3664 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=145110 $Y=12870 $D=28
M3208 3667 3666 3665 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=145670 $Y=12870 $D=28
M3209 3677 3663 3667 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=146230 $Y=13110 $D=28
M3210 VSS 3669 3677 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=146550 $Y=13110 $D=28
M3211 3678 584 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=146990 $Y=13090 $D=28
M3212 3669 3667 3678 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=147310 $Y=13090 $D=28
M3213 3668 3669 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=147630 $Y=12390 $D=28
M3214 VSS 3668 3661 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=148530 $Y=13070 $D=28
M3215 result[19] 3669 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=149030 $Y=13070 $D=28
M3216 3686 3679 3680 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=150060 $Y=13090 $D=28
M3217 3688 623 3686 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=150380 $Y=13090 $D=28
M3218 VSS 638 3688 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=150700 $Y=13090 $D=28
M3219 VSS clk 3679 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=151680 $Y=12840 $D=28
M3220 3682 3679 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=152190 $Y=12940 $D=28
M3221 3690 3682 3680 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=153210 $Y=13010 $D=28
M3222 3691 3681 3690 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=153530 $Y=13010 $D=28
M3223 VSS 638 3691 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=153850 $Y=13010 $D=28
M3224 3681 3680 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=154310 $Y=12870 $D=28
M3225 3683 3682 3681 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=154870 $Y=12870 $D=28
M3226 3693 3679 3683 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=155430 $Y=13110 $D=28
M3227 VSS 3685 3693 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=155750 $Y=13110 $D=28
M3228 3694 638 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=156190 $Y=13090 $D=28
M3229 3685 3683 3694 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=156510 $Y=13090 $D=28
M3230 3684 3685 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=156830 $Y=12390 $D=28
M3231 VSS 3684 3662 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=157730 $Y=13070 $D=28
M3232 result[20] 3685 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=158230 $Y=13070 $D=28
M3233 3704 3697 3698 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=149260 $Y=27490 $D=28
M3234 3706 612 3704 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=149580 $Y=27490 $D=28
M3235 VSS 662 3706 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=149900 $Y=27490 $D=28
M3236 VSS clk 3697 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=150880 $Y=27240 $D=28
M3237 3700 3697 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=151390 $Y=27340 $D=28
M3238 3708 3700 3698 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=152410 $Y=27410 $D=28
M3239 3709 3699 3708 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=152730 $Y=27410 $D=28
M3240 VSS 662 3709 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=153050 $Y=27410 $D=28
M3241 3699 3698 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=153510 $Y=27270 $D=28
M3242 3701 3700 3699 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=154070 $Y=27270 $D=28
M3243 3711 3697 3701 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=154630 $Y=27510 $D=28
M3244 VSS 3703 3711 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=154950 $Y=27510 $D=28
M3245 3712 662 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=155390 $Y=27490 $D=28
M3246 3703 3701 3712 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=155710 $Y=27490 $D=28
M3247 3702 3703 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=156030 $Y=26790 $D=28
M3248 VSS 3702 3695 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=156930 $Y=27470 $D=28
M3249 result[25] 3703 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=157430 $Y=27470 $D=28
M3250 3720 3713 3714 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=158460 $Y=27490 $D=28
M3251 3722 656 3720 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=158780 $Y=27490 $D=28
M3252 VSS 641 3722 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=159100 $Y=27490 $D=28
M3253 VSS clk 3713 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=160080 $Y=27240 $D=28
M3254 3716 3713 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=160590 $Y=27340 $D=28
M3255 3724 3716 3714 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=161610 $Y=27410 $D=28
M3256 3725 3715 3724 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=161930 $Y=27410 $D=28
M3257 VSS 641 3725 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=162250 $Y=27410 $D=28
M3258 3715 3714 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=162710 $Y=27270 $D=28
M3259 3717 3716 3715 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=163270 $Y=27270 $D=28
M3260 3727 3713 3717 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=163830 $Y=27510 $D=28
M3261 VSS 3719 3727 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.5766e-14 as=2e-14 pd=5.29787e-07 ps=4e-07 nrd=1.89415 nrs=0.5 sa=6.6e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=164150 $Y=27510 $D=28
M3262 3728 641 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.2e-14 as=8.33426e-14 pd=4.2e-07 ps=5.82766e-07 nrd=0.454545 nrs=1.72195 sa=1.02182e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=164590 $Y=27490 $D=28
M3263 3719 3717 3728 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=2.2e-14 pd=1.28e-06 ps=4.2e-07 nrd=1.98347 nrs=0.454545 sa=1.34182e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=164910 $Y=27490 $D=28
M3264 3718 3719 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.5766e-14 pd=1.28e-06 ps=5.29787e-07 nrd=2.36 nrs=1.89415 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=165230 $Y=26790 $D=28
M3265 VSS 3718 3696 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02758e-13 as=9.76e-14 pd=1.02947e-06 ps=1.28e-06 nrd=1.78399 nrs=1.69444 sa=3.6e-07 sb=8.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=166130 $Y=27470 $D=28
M3266 result[26] 3719 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.76e-14 as=1.02758e-13 pd=1.28e-06 ps=1.02947e-06 nrd=1.69444 nrs=1.78399 sa=8.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=166630 $Y=27470 $D=28
M3267 VSS 228 3729 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.85556e-14 as=9.44e-14 pd=5.81481e-07 ps=1.28e-06 nrd=1.71389 nrs=2.36 sa=3.6e-07 sb=1.18e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=61760 $Y=53950 $D=28
M3268 3730 241 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.05667e-13 pd=8e-07 ps=1.74444e-06 nrd=0.166667 nrs=0.571296 sa=5.29667e-07 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=62300 $Y=53950 $D=28
M3269 221 3729 3730 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=8.49667e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=62620 $Y=53950 $D=28
M3270 VSS 437 3731 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.85556e-14 as=9.44e-14 pd=5.81481e-07 ps=1.28e-06 nrd=1.71389 nrs=2.36 sa=3.6e-07 sb=1.18e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=112560 $Y=56250 $D=28
M3271 3732 430 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.05667e-13 pd=8e-07 ps=1.74444e-06 nrd=0.166667 nrs=0.571296 sa=5.29667e-07 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=113100 $Y=55850 $D=28
M3272 412 3731 3732 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=8.49667e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=113420 $Y=55850 $D=28
M3273 VSS 562 3733 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.85556e-14 as=9.44e-14 pd=5.81481e-07 ps=1.28e-06 nrd=1.71389 nrs=2.36 sa=3.6e-07 sb=1.18e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=138160 $Y=68350 $D=28
M3274 3734 539 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.05667e-13 pd=8e-07 ps=1.74444e-06 nrd=0.166667 nrs=0.571296 sa=5.29667e-07 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=138700 $Y=68350 $D=28
M3275 913 3733 3734 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=8.49667e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=139020 $Y=68350 $D=28
M3276 VSS 559 3735 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.85556e-14 as=9.44e-14 pd=5.81481e-07 ps=1.28e-06 nrd=1.71389 nrs=2.36 sa=3.6e-07 sb=1.18e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=138560 $Y=61150 $D=28
M3277 3736 549 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.05667e-13 pd=8e-07 ps=1.74444e-06 nrd=0.166667 nrs=0.571296 sa=5.29667e-07 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=139100 $Y=61150 $D=28
M3278 553 3735 3736 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=8.49667e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=139420 $Y=61150 $D=28
M3279 VSS 575 3737 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.85556e-14 as=9.44e-14 pd=5.81481e-07 ps=1.28e-06 nrd=1.71389 nrs=2.36 sa=3.6e-07 sb=1.18e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=143760 $Y=61150 $D=28
M3280 3738 560 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6e-14 as=2.05667e-13 pd=8e-07 ps=1.74444e-06 nrd=0.166667 nrs=0.571296 sa=5.29667e-07 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=144300 $Y=61150 $D=28
M3281 567 3737 3738 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=6e-14 pd=1.84e-06 ps=8e-07 nrd=0.533333 nrs=0.166667 sa=8.49667e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=144620 $Y=61150 $D=28
M3282 87 82 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.72419e-13 as=2.944e-13 pd=1.38541e-06 ps=2.48e-06 nrd=0.203708 nrs=0.347826 sa=3.2e-07 sb=7.19348e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=26810 $Y=55590 $D=28
M3283 VSS 82 87 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.46181e-13 pd=2.2e-06 ps=1.17459e-06 nrd=0.410256 nrs=0.240271 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=27290 $Y=55730 $D=28
M3284 148 97 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.72419e-13 as=2.944e-13 pd=1.38541e-06 ps=2.48e-06 nrd=0.203708 nrs=0.347826 sa=3.2e-07 sb=7.19348e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=40810 $Y=25090 $D=28
M3285 VSS 97 148 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.46181e-13 pd=2.2e-06 ps=1.17459e-06 nrd=0.410256 nrs=0.240271 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=41290 $Y=25090 $D=28
M3286 411 402 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.72419e-13 as=2.944e-13 pd=1.38541e-06 ps=2.48e-06 nrd=0.203708 nrs=0.347826 sa=3.2e-07 sb=7.19348e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=108010 $Y=75490 $D=28
M3287 VSS 402 411 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.46181e-13 pd=2.2e-06 ps=1.17459e-06 nrd=0.410256 nrs=0.240271 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=108490 $Y=75490 $D=28
M3288 435 404 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.72419e-13 as=2.944e-13 pd=1.38541e-06 ps=2.48e-06 nrd=0.203708 nrs=0.347826 sa=3.2e-07 sb=7.19348e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=110810 $Y=69990 $D=28
M3289 VSS 404 435 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.46181e-13 pd=2.2e-06 ps=1.17459e-06 nrd=0.410256 nrs=0.240271 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=111290 $Y=70130 $D=28
M3290 499 523 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.72419e-13 as=2.944e-13 pd=1.38541e-06 ps=2.48e-06 nrd=0.203708 nrs=0.347826 sa=3.2e-07 sb=7.19348e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=133210 $Y=39490 $D=28
M3291 VSS 523 499 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.46181e-13 pd=2.2e-06 ps=1.17459e-06 nrd=0.410256 nrs=0.240271 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=133690 $Y=39490 $D=28
M3292 849 503 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.72419e-13 as=2.944e-13 pd=1.38541e-06 ps=2.48e-06 nrd=0.203708 nrs=0.347826 sa=3.2e-07 sb=7.19348e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=133610 $Y=68290 $D=28
M3293 VSS 503 849 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.46181e-13 pd=2.2e-06 ps=1.17459e-06 nrd=0.410256 nrs=0.240271 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=134090 $Y=68290 $D=28
M3294 VSS 59 3739 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=2.944e-13 pd=1.61247e-06 ps=2.48e-06 nrd=0.200561 nrs=0.347826 sa=3.2e-07 sb=1.50261e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=20450 $Y=53890 $D=28
M3295 3739 63 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20972e-13 as=1.21781e-13 pd=1.06937e-06 ps=1.15677e-06 nrd=0.277714 nrs=0.27957 sa=7.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=20890 $Y=53890 $D=28
M3296 VSS 63 3739 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=1.68628e-13 pd=1.61247e-06 ps=1.49063e-06 nrd=0.200561 nrs=0.199229 sa=9.46087e-07 sb=1.48696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=21370 $Y=53890 $D=28
M3297 3739 59 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=1.21781e-13 pd=1.02e-06 ps=1.15677e-06 nrd=0.272727 nrs=0.27957 sa=1.68e-06 sb=1.95152e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=21810 $Y=53890 $D=28
M3298 VSS 59 3739 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3299e-13 as=1.188e-13 pd=1.34475e-06 ps=1.02e-06 nrd=0.305303 nrs=0.272727 sa=2e-06 sb=1.92242e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=22290 $Y=53890 $D=28
M3299 3739 63 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22368e-13 as=1.3299e-13 pd=1.08811e-06 ps=1.34475e-06 nrd=0.280917 nrs=0.305303 sa=2e-06 sb=1.6703e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=22730 $Y=53890 $D=28
M3300 803 75 3739 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.52032e-13 pd=1.18e-06 ps=1.35189e-06 nrd=0.219512 nrs=0.226104 sa=1.56098e-06 sb=1.28e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=23210 $Y=53930 $D=28
M3301 3739 75 803 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.67805e-06 sb=8e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=23690 $Y=53930 $D=28
M3302 803 75 3739 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.79512e-06 sb=3.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=24170 $Y=53930 $D=28
M3303 VSS 142 3743 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=2.944e-13 pd=1.61247e-06 ps=2.48e-06 nrd=0.200561 nrs=0.347826 sa=3.2e-07 sb=1.50261e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1e-15 $X=29650 $Y=41190 $D=28
M3304 3743 84 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20972e-13 as=1.21781e-13 pd=1.06937e-06 ps=1.15677e-06 nrd=0.277714 nrs=0.27957 sa=7.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=30090 $Y=41450 $D=28
M3305 VSS 84 3743 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=1.68628e-13 pd=1.61247e-06 ps=1.49063e-06 nrd=0.200561 nrs=0.199229 sa=9.46087e-07 sb=1.48696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=1.2e-14 $X=30570 $Y=41190 $D=28
M3306 3743 142 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=1.21781e-13 pd=1.02e-06 ps=1.15677e-06 nrd=0.272727 nrs=0.27957 sa=1.68e-06 sb=1.95152e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=31010 $Y=41450 $D=28
M3307 VSS 142 3743 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3299e-13 as=1.188e-13 pd=1.34475e-06 ps=1.02e-06 nrd=0.305303 nrs=0.272727 sa=2e-06 sb=1.92242e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=31490 $Y=41450 $D=28
M3308 3743 84 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22368e-13 as=1.3299e-13 pd=1.08811e-06 ps=1.34475e-06 nrd=0.280917 nrs=0.305303 sa=2e-06 sb=1.6703e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=31930 $Y=41450 $D=28
M3309 103 108 3743 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.52032e-13 pd=1.18e-06 ps=1.35189e-06 nrd=0.219512 nrs=0.226104 sa=1.56098e-06 sb=1.28e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=32410 $Y=41250 $D=28
M3310 3743 108 103 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.67805e-06 sb=8e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=32890 $Y=41250 $D=28
M3311 103 108 3743 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.79512e-06 sb=3.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=33370 $Y=41250 $D=28
M3312 VSS 119 3747 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=2.944e-13 pd=1.61247e-06 ps=2.48e-06 nrd=0.200561 nrs=0.347826 sa=3.2e-07 sb=1.50261e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=30050 $Y=19590 $D=28
M3313 3747 118 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20972e-13 as=1.21781e-13 pd=1.06937e-06 ps=1.15677e-06 nrd=0.277714 nrs=0.27957 sa=7.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=30490 $Y=19850 $D=28
M3314 VSS 118 3747 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=1.68628e-13 pd=1.61247e-06 ps=1.49063e-06 nrd=0.200561 nrs=0.199229 sa=9.46087e-07 sb=1.48696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=30970 $Y=19590 $D=28
M3315 3747 119 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=1.21781e-13 pd=1.02e-06 ps=1.15677e-06 nrd=0.272727 nrs=0.27957 sa=1.68e-06 sb=1.95152e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=31410 $Y=19850 $D=28
M3316 VSS 119 3747 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3299e-13 as=1.188e-13 pd=1.34475e-06 ps=1.02e-06 nrd=0.305303 nrs=0.272727 sa=2e-06 sb=1.92242e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=31890 $Y=19850 $D=28
M3317 3747 118 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22368e-13 as=1.3299e-13 pd=1.08811e-06 ps=1.34475e-06 nrd=0.280917 nrs=0.305303 sa=2e-06 sb=1.6703e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=32330 $Y=19850 $D=28
M3318 15 132 3747 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.52032e-13 pd=1.18e-06 ps=1.35189e-06 nrd=0.219512 nrs=0.226104 sa=1.56098e-06 sb=1.28e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=32810 $Y=19650 $D=28
M3319 3747 132 15 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.67805e-06 sb=8e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=33290 $Y=19650 $D=28
M3320 15 132 3747 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.79512e-06 sb=3.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=33770 $Y=19650 $D=28
M3321 VSS 143 3751 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=2.944e-13 pd=1.61247e-06 ps=2.48e-06 nrd=0.200561 nrs=0.347826 sa=3.2e-07 sb=1.50261e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=41250 $Y=17890 $D=28
M3322 3751 177 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20972e-13 as=1.21781e-13 pd=1.06937e-06 ps=1.15677e-06 nrd=0.277714 nrs=0.27957 sa=7.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=41690 $Y=17890 $D=28
M3323 VSS 177 3751 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=1.68628e-13 pd=1.61247e-06 ps=1.49063e-06 nrd=0.200561 nrs=0.199229 sa=9.46087e-07 sb=1.48696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=42170 $Y=17890 $D=28
M3324 3751 143 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=1.21781e-13 pd=1.02e-06 ps=1.15677e-06 nrd=0.272727 nrs=0.27957 sa=1.68e-06 sb=1.95152e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=42610 $Y=17890 $D=28
M3325 VSS 143 3751 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3299e-13 as=1.188e-13 pd=1.34475e-06 ps=1.02e-06 nrd=0.305303 nrs=0.272727 sa=2e-06 sb=1.92242e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=43090 $Y=17890 $D=28
M3326 3751 177 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22368e-13 as=1.3299e-13 pd=1.08811e-06 ps=1.34475e-06 nrd=0.280917 nrs=0.305303 sa=2e-06 sb=1.6703e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=43530 $Y=17890 $D=28
M3327 167 169 3751 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.52032e-13 pd=1.18e-06 ps=1.35189e-06 nrd=0.219512 nrs=0.226104 sa=1.56098e-06 sb=1.28e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=44010 $Y=17930 $D=28
M3328 3751 169 167 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.67805e-06 sb=8e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=44490 $Y=17930 $D=28
M3329 167 169 3751 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.79512e-06 sb=3.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=44970 $Y=17930 $D=28
M3330 VSS 358 3755 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=2.944e-13 pd=1.61247e-06 ps=2.48e-06 nrd=0.200561 nrs=0.347826 sa=3.2e-07 sb=1.50261e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=95650 $Y=75490 $D=28
M3331 3755 353 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20972e-13 as=1.21781e-13 pd=1.06937e-06 ps=1.15677e-06 nrd=0.277714 nrs=0.27957 sa=7.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=96090 $Y=75490 $D=28
M3332 VSS 353 3755 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=1.68628e-13 pd=1.61247e-06 ps=1.49063e-06 nrd=0.200561 nrs=0.199229 sa=9.46087e-07 sb=1.48696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=96570 $Y=75490 $D=28
M3333 3755 358 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=1.21781e-13 pd=1.02e-06 ps=1.15677e-06 nrd=0.272727 nrs=0.27957 sa=1.68e-06 sb=1.95152e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=97010 $Y=75490 $D=28
M3334 VSS 358 3755 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3299e-13 as=1.188e-13 pd=1.34475e-06 ps=1.02e-06 nrd=0.305303 nrs=0.272727 sa=2e-06 sb=1.92242e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=97490 $Y=75490 $D=28
M3335 3755 353 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22368e-13 as=1.3299e-13 pd=1.08811e-06 ps=1.34475e-06 nrd=0.280917 nrs=0.305303 sa=2e-06 sb=1.6703e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=97930 $Y=75490 $D=28
M3336 404 361 3755 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.52032e-13 pd=1.18e-06 ps=1.35189e-06 nrd=0.219512 nrs=0.226104 sa=1.56098e-06 sb=1.28e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=98410 $Y=75530 $D=28
M3337 3755 361 404 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.67805e-06 sb=8e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=98890 $Y=75530 $D=28
M3338 404 361 3755 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.79512e-06 sb=3.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=99370 $Y=75530 $D=28
M3339 VSS 496 3759 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=2.944e-13 pd=1.61247e-06 ps=2.48e-06 nrd=0.200561 nrs=0.347826 sa=3.2e-07 sb=1.50261e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=122050 $Y=69990 $D=28
M3340 3759 402 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20972e-13 as=1.21781e-13 pd=1.06937e-06 ps=1.15677e-06 nrd=0.277714 nrs=0.27957 sa=7.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=122490 $Y=70250 $D=28
M3341 VSS 402 3759 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=1.68628e-13 pd=1.61247e-06 ps=1.49063e-06 nrd=0.200561 nrs=0.199229 sa=9.46087e-07 sb=1.48696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=122970 $Y=69990 $D=28
M3342 3759 496 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=1.21781e-13 pd=1.02e-06 ps=1.15677e-06 nrd=0.272727 nrs=0.27957 sa=1.68e-06 sb=1.95152e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=123410 $Y=70250 $D=28
M3343 VSS 496 3759 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3299e-13 as=1.188e-13 pd=1.34475e-06 ps=1.02e-06 nrd=0.305303 nrs=0.272727 sa=2e-06 sb=1.92242e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=123890 $Y=70250 $D=28
M3344 3759 402 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22368e-13 as=1.3299e-13 pd=1.08811e-06 ps=1.34475e-06 nrd=0.280917 nrs=0.305303 sa=2e-06 sb=1.6703e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=124330 $Y=70250 $D=28
M3345 503 842 3759 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.52032e-13 pd=1.18e-06 ps=1.35189e-06 nrd=0.219512 nrs=0.226104 sa=1.56098e-06 sb=1.28e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=124810 $Y=70050 $D=28
M3346 3759 842 503 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.67805e-06 sb=8e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=125290 $Y=70050 $D=28
M3347 503 842 3759 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.79512e-06 sb=3.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=125770 $Y=70050 $D=28
M3348 VSS 476 3763 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=2.944e-13 pd=1.61247e-06 ps=2.48e-06 nrd=0.200561 nrs=0.347826 sa=3.2e-07 sb=1.50261e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=126850 $Y=68290 $D=28
M3349 3763 846 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20972e-13 as=1.21781e-13 pd=1.06937e-06 ps=1.15677e-06 nrd=0.277714 nrs=0.27957 sa=7.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=127290 $Y=68290 $D=28
M3350 VSS 846 3763 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=1.68628e-13 pd=1.61247e-06 ps=1.49063e-06 nrd=0.200561 nrs=0.199229 sa=9.46087e-07 sb=1.48696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=127770 $Y=68290 $D=28
M3351 3763 476 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=1.21781e-13 pd=1.02e-06 ps=1.15677e-06 nrd=0.272727 nrs=0.27957 sa=1.68e-06 sb=1.95152e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=128210 $Y=68290 $D=28
M3352 VSS 476 3763 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3299e-13 as=1.188e-13 pd=1.34475e-06 ps=1.02e-06 nrd=0.305303 nrs=0.272727 sa=2e-06 sb=1.92242e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=128690 $Y=68290 $D=28
M3353 3763 846 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22368e-13 as=1.3299e-13 pd=1.08811e-06 ps=1.34475e-06 nrd=0.280917 nrs=0.305303 sa=2e-06 sb=1.6703e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=129130 $Y=68290 $D=28
M3354 482 495 3763 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.52032e-13 pd=1.18e-06 ps=1.35189e-06 nrd=0.219512 nrs=0.226104 sa=1.56098e-06 sb=1.28e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=129610 $Y=68330 $D=28
M3355 3763 495 482 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.67805e-06 sb=8e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=130090 $Y=68330 $D=28
M3356 482 495 3763 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.79512e-06 sb=3.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=130570 $Y=68330 $D=28
M3357 VSS 502 3767 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=2.944e-13 pd=1.61247e-06 ps=2.48e-06 nrd=0.200561 nrs=0.347826 sa=3.2e-07 sb=1.50261e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=132450 $Y=46690 $D=28
M3358 3767 512 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20972e-13 as=1.21781e-13 pd=1.06937e-06 ps=1.15677e-06 nrd=0.277714 nrs=0.27957 sa=7.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=132890 $Y=46690 $D=28
M3359 VSS 512 3767 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69755e-13 as=1.68628e-13 pd=1.61247e-06 ps=1.49063e-06 nrd=0.200561 nrs=0.199229 sa=9.46087e-07 sb=1.48696e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=133370 $Y=46690 $D=28
M3360 3767 502 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=1.21781e-13 pd=1.02e-06 ps=1.15677e-06 nrd=0.272727 nrs=0.27957 sa=1.68e-06 sb=1.95152e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=133810 $Y=46690 $D=28
M3361 VSS 502 3767 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3299e-13 as=1.188e-13 pd=1.34475e-06 ps=1.02e-06 nrd=0.305303 nrs=0.272727 sa=2e-06 sb=1.92242e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=134290 $Y=46690 $D=28
M3362 3767 512 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22368e-13 as=1.3299e-13 pd=1.08811e-06 ps=1.34475e-06 nrd=0.280917 nrs=0.305303 sa=2e-06 sb=1.6703e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=134730 $Y=46690 $D=28
M3363 598 532 3767 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.52032e-13 pd=1.18e-06 ps=1.35189e-06 nrd=0.219512 nrs=0.226104 sa=1.56098e-06 sb=1.28e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=135210 $Y=46730 $D=28
M3364 3767 532 598 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.67805e-06 sb=8e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=135690 $Y=46730 $D=28
M3365 598 532 3767 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.79512e-06 sb=3.2e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=136170 $Y=46730 $D=28
M3366 78 112 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.67043e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=33210 $Y=33990 $D=28
M3367 VSS 112 78 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8e-07 sb=1.19043e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=33690 $Y=33990 $D=28
M3368 78 112 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.68628e-13 as=2.08475e-13 pd=1.49063e-06 ps=1.41472e-06 nrd=0.199229 nrs=0.246308 sa=1.36e-06 sb=6.30435e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=34250 $Y=33990 $D=28
M3369 VSS 112 78 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.112e-13 as=1.20972e-13 pd=1.96e-06 ps=1.06937e-06 nrd=0.484848 nrs=0.277714 sa=1.84e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=34730 $Y=34250 $D=28
M3370 123 112 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.67043e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=6e-15 $X=34410 $Y=41190 $D=28
M3371 VSS 112 123 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8e-07 sb=1.19043e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=6e-15 $X=34890 $Y=41190 $D=28
M3372 123 112 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.68628e-13 as=2.08475e-13 pd=1.49063e-06 ps=1.41472e-06 nrd=0.199229 nrs=0.246308 sa=1.36e-06 sb=6.30435e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=6e-15 $X=35450 $Y=41190 $D=28
M3373 VSS 112 123 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.112e-13 as=1.20972e-13 pd=1.96e-06 ps=1.06937e-06 nrd=0.484848 nrs=0.277714 sa=1.84e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=35930 $Y=41450 $D=28
M3374 278 236 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.67043e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=58410 $Y=32290 $D=28
M3375 VSS 236 278 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8e-07 sb=1.19043e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=58890 $Y=32290 $D=28
M3376 278 236 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.68628e-13 as=2.08475e-13 pd=1.49063e-06 ps=1.41472e-06 nrd=0.199229 nrs=0.246308 sa=1.36e-06 sb=6.30435e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=59450 $Y=32290 $D=28
M3377 VSS 236 278 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.112e-13 as=1.20972e-13 pd=1.96e-06 ps=1.06937e-06 nrd=0.484848 nrs=0.277714 sa=1.84e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=59930 $Y=32290 $D=28
M3378 231 263 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.67043e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=61210 $Y=32290 $D=28
M3379 VSS 263 231 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8e-07 sb=1.19043e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=61690 $Y=32290 $D=28
M3380 231 263 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.68628e-13 as=2.08475e-13 pd=1.49063e-06 ps=1.41472e-06 nrd=0.199229 nrs=0.246308 sa=1.36e-06 sb=6.30435e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=62250 $Y=32290 $D=28
M3381 VSS 263 231 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.112e-13 as=1.20972e-13 pd=1.96e-06 ps=1.06937e-06 nrd=0.484848 nrs=0.277714 sa=1.84e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=62730 $Y=32290 $D=28
M3382 301 284 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.67043e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=75610 $Y=39490 $D=28
M3383 VSS 284 301 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8e-07 sb=1.19043e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=76090 $Y=39490 $D=28
M3384 301 284 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.68628e-13 as=2.08475e-13 pd=1.49063e-06 ps=1.41472e-06 nrd=0.199229 nrs=0.246308 sa=1.36e-06 sb=6.30435e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=76650 $Y=39490 $D=28
M3385 VSS 284 301 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.112e-13 as=1.20972e-13 pd=1.96e-06 ps=1.06937e-06 nrd=0.484848 nrs=0.277714 sa=1.84e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=77130 $Y=39490 $D=28
M3386 523 503 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.67043e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=131210 $Y=62790 $D=28
M3387 VSS 503 523 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=8e-07 sb=1.19043e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=131690 $Y=62790 $D=28
M3388 523 503 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.68628e-13 as=2.08475e-13 pd=1.49063e-06 ps=1.41472e-06 nrd=0.199229 nrs=0.246308 sa=1.36e-06 sb=6.30435e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=132250 $Y=62790 $D=28
M3389 VSS 503 523 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.112e-13 as=1.20972e-13 pd=1.96e-06 ps=1.06937e-06 nrd=0.484848 nrs=0.277714 sa=1.84e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=132730 $Y=63050 $D=28
M3390 3773 49 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=18430 $Y=27160 $D=28
M3391 VSS 49 3773 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=18910 $Y=27160 $D=28
M3392 3772 3773 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=19350 $Y=27160 $D=28
M3393 VSS 3773 3772 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=19830 $Y=27160 $D=28
M3394 3771 78 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=20270 $Y=27110 $D=28
M3395 3772 78 57 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=21230 $Y=27000 $D=28
M3396 57 78 3772 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=21710 $Y=27000 $D=28
M3397 3773 3771 57 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=22190 $Y=27000 $D=28
M3398 57 3771 3773 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=22670 $Y=27000 $D=28
M3399 3776 127 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=25630 $Y=34360 $D=28
M3400 VSS 127 3776 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=26110 $Y=34360 $D=28
M3401 3775 3776 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=26550 $Y=34360 $D=28
M3402 VSS 3776 3775 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=27030 $Y=34360 $D=28
M3403 3774 123 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=27470 $Y=34310 $D=28
M3404 3775 123 107 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=28430 $Y=34200 $D=28
M3405 107 123 3775 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=28910 $Y=34200 $D=28
M3406 3776 3774 107 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=29390 $Y=34200 $D=28
M3407 107 3774 3776 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=29870 $Y=34200 $D=28
M3408 3779 136 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=32030 $Y=46690 $D=28
M3409 VSS 136 3779 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=32510 $Y=46690 $D=28
M3410 3778 3779 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=32950 $Y=46690 $D=28
M3411 VSS 3779 3778 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=33430 $Y=46690 $D=28
M3412 3777 123 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=33870 $Y=46850 $D=28
M3413 3778 123 131 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=34830 $Y=46850 $D=28
M3414 131 123 3778 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=35310 $Y=46850 $D=28
M3415 3779 3777 131 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=35790 $Y=46850 $D=28
M3416 131 3777 3779 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=36270 $Y=46850 $D=28
M3417 3782 141 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=34030 $Y=32290 $D=28
M3418 VSS 141 3782 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=34510 $Y=32290 $D=28
M3419 3781 3782 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=34950 $Y=32290 $D=28
M3420 VSS 3782 3781 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=35430 $Y=32290 $D=28
M3421 3780 78 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=35870 $Y=32450 $D=28
M3422 3781 78 142 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=36830 $Y=32450 $D=28
M3423 142 78 3781 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=37310 $Y=32450 $D=28
M3424 3782 3780 142 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=37790 $Y=32450 $D=28
M3425 142 3780 3782 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=38270 $Y=32450 $D=28
M3426 3785 127 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=36030 $Y=34360 $D=28
M3427 VSS 127 3785 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=36510 $Y=34360 $D=28
M3428 3784 3785 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=36950 $Y=34360 $D=28
M3429 VSS 3785 3784 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=37430 $Y=34360 $D=28
M3430 3783 123 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=37870 $Y=34310 $D=28
M3431 3784 123 893 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=38830 $Y=34200 $D=28
M3432 893 123 3784 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=39310 $Y=34200 $D=28
M3433 3785 3783 893 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=39790 $Y=34200 $D=28
M3434 893 3783 3785 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=40270 $Y=34200 $D=28
M3435 3788 157 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=40030 $Y=41560 $D=28
M3436 VSS 157 3788 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=40510 $Y=41560 $D=28
M3437 3787 3788 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=40950 $Y=41560 $D=28
M3438 VSS 3788 3787 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=41430 $Y=41560 $D=28
M3439 3786 163 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=41870 $Y=41510 $D=28
M3440 3787 163 166 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=42830 $Y=41400 $D=28
M3441 166 163 3787 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=43310 $Y=41400 $D=28
M3442 3788 3786 166 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=43790 $Y=41400 $D=28
M3443 166 3786 3788 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=44270 $Y=41400 $D=28
M3444 3791 157 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=40430 $Y=53890 $D=28
M3445 VSS 157 3791 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=40910 $Y=53890 $D=28
M3446 3790 3791 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=41350 $Y=53890 $D=28
M3447 VSS 3791 3790 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=41830 $Y=53890 $D=28
M3448 3789 78 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=42270 $Y=54050 $D=28
M3449 3790 78 174 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=43230 $Y=54050 $D=28
M3450 174 78 3790 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=43710 $Y=54050 $D=28
M3451 3791 3789 174 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=44190 $Y=54050 $D=28
M3452 174 3789 3791 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=44670 $Y=54050 $D=28
M3453 3794 78 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=43630 $Y=55960 $D=28
M3454 VSS 78 3794 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=44110 $Y=55960 $D=28
M3455 3793 3794 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=44550 $Y=55960 $D=28
M3456 VSS 3794 3793 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=45030 $Y=55960 $D=28
M3457 3792 186 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=45470 $Y=55910 $D=28
M3458 3793 186 181 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=46430 $Y=55800 $D=28
M3459 181 186 3793 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=46910 $Y=55800 $D=28
M3460 3794 3792 181 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=47390 $Y=55800 $D=28
M3461 181 3792 3794 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=47870 $Y=55800 $D=28
M3462 3797 171 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=45630 $Y=53890 $D=28
M3463 VSS 171 3797 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=46110 $Y=53890 $D=28
M3464 3796 3797 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=46550 $Y=53890 $D=28
M3465 VSS 3797 3796 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=47030 $Y=53890 $D=28
M3466 3795 78 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=47470 $Y=54050 $D=28
M3467 3796 78 179 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=48430 $Y=54050 $D=28
M3468 179 78 3796 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=48910 $Y=54050 $D=28
M3469 3797 3795 179 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=49390 $Y=54050 $D=28
M3470 179 3795 3797 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=49870 $Y=54050 $D=28
M3471 3800 240 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=74830 $Y=27160 $D=28
M3472 VSS 240 3800 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=75310 $Y=27160 $D=28
M3473 3799 3800 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=75750 $Y=27160 $D=28
M3474 VSS 3800 3799 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=76230 $Y=27160 $D=28
M3475 3798 287 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=76670 $Y=27110 $D=28
M3476 3799 287 280 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=77630 $Y=27000 $D=28
M3477 280 287 3799 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=78110 $Y=27000 $D=28
M3478 3800 3798 280 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=78590 $Y=27000 $D=28
M3479 280 3798 3800 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=79070 $Y=27000 $D=28
M3480 3803 240 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=74830 $Y=32290 $D=28
M3481 VSS 240 3803 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=75310 $Y=32290 $D=28
M3482 3802 3803 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=75750 $Y=32290 $D=28
M3483 VSS 3803 3802 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=76230 $Y=32290 $D=28
M3484 3801 254 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=76670 $Y=32450 $D=28
M3485 3802 254 293 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=77630 $Y=32450 $D=28
M3486 293 254 3802 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=78110 $Y=32450 $D=28
M3487 3803 3801 293 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=78590 $Y=32450 $D=28
M3488 293 3801 3803 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=79070 $Y=32450 $D=28
M3489 3806 157 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=79230 $Y=46690 $D=28
M3490 VSS 157 3806 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=79710 $Y=46690 $D=28
M3491 3805 3806 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=80150 $Y=46690 $D=28
M3492 VSS 3806 3805 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=80630 $Y=46690 $D=28
M3493 3804 307 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=81070 $Y=46850 $D=28
M3494 3805 307 319 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=82030 $Y=46850 $D=28
M3495 319 307 3805 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=82510 $Y=46850 $D=28
M3496 3806 3804 319 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=82990 $Y=46850 $D=28
M3497 319 3804 3806 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=83470 $Y=46850 $D=28
M3498 3809 186 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=80430 $Y=55960 $D=28
M3499 VSS 186 3809 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=80910 $Y=55960 $D=28
M3500 3808 3809 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=81350 $Y=55960 $D=28
M3501 VSS 3809 3808 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=81830 $Y=55960 $D=28
M3502 3807 307 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=82270 $Y=55910 $D=28
M3503 3808 307 314 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=83230 $Y=55800 $D=28
M3504 314 307 3808 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=83710 $Y=55800 $D=28
M3505 3809 3807 314 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=84190 $Y=55800 $D=28
M3506 314 3807 3809 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=84670 $Y=55800 $D=28
M3507 3812 354 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=84030 $Y=34360 $D=28
M3508 VSS 354 3812 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=84510 $Y=34360 $D=28
M3509 3811 3812 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=84950 $Y=34360 $D=28
M3510 VSS 3812 3811 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=85430 $Y=34360 $D=28
M3511 3810 192 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=85870 $Y=34310 $D=28
M3512 3811 192 328 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=86830 $Y=34200 $D=28
M3513 328 192 3811 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=87310 $Y=34200 $D=28
M3514 3812 3810 328 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=87790 $Y=34200 $D=28
M3515 328 3810 3812 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=88270 $Y=34200 $D=28
M3516 3815 171 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=84430 $Y=46690 $D=28
M3517 VSS 171 3815 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=84910 $Y=46690 $D=28
M3518 3814 3815 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=85350 $Y=46690 $D=28
M3519 VSS 3815 3814 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=85830 $Y=46690 $D=28
M3520 3813 307 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=86270 $Y=46850 $D=28
M3521 3814 307 327 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=87230 $Y=46850 $D=28
M3522 327 307 3814 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=87710 $Y=46850 $D=28
M3523 3815 3813 327 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=88190 $Y=46850 $D=28
M3524 327 3813 3815 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=88670 $Y=46850 $D=28
M3525 3818 176 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=88430 $Y=39490 $D=28
M3526 VSS 176 3818 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=88910 $Y=39490 $D=28
M3527 3817 3818 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=89350 $Y=39490 $D=28
M3528 VSS 3818 3817 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=89830 $Y=39490 $D=28
M3529 3816 354 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=90270 $Y=39650 $D=28
M3530 3817 354 343 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=91230 $Y=39650 $D=28
M3531 343 354 3817 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=91710 $Y=39650 $D=28
M3532 3818 3816 343 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=92190 $Y=39650 $D=28
M3533 343 3816 3818 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=92670 $Y=39650 $D=28
M3534 3821 538 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=104830 $Y=48760 $D=28
M3535 VSS 538 3821 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=105310 $Y=48760 $D=28
M3536 3820 3821 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=105750 $Y=48760 $D=28
M3537 VSS 3821 3820 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=106230 $Y=48760 $D=28
M3538 3819 395 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=106670 $Y=48710 $D=28
M3539 3820 395 406 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=107630 $Y=48600 $D=28
M3540 406 395 3820 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=108110 $Y=48600 $D=28
M3541 3821 3819 406 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=108590 $Y=48600 $D=28
M3542 406 3819 3821 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=109070 $Y=48600 $D=28
M3543 3824 520 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.87e-13 pd=9.1e-07 ps=1.78e-06 nrd=0.327273 nrs=0.618182 sa=3.4e-07 sb=1.88364e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=127630 $Y=53890 $D=28
M3544 VSS 520 3824 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24348e-13 as=9.9e-14 pd=1.29928e-06 ps=9.1e-07 nrd=0.411067 nrs=0.327273 sa=8.2e-07 sb=1.51709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=128110 $Y=53890 $D=28
M3545 3823 3824 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.24348e-13 pd=9.1e-07 ps=1.29928e-06 nrd=0.327273 nrs=0.411067 sa=1.26e-06 sb=1.07709e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=128550 $Y=53890 $D=28
M3546 VSS 3824 3823 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28535e-13 as=9.9e-14 pd=1.41181e-06 ps=9.1e-07 nrd=0.424911 nrs=0.327273 sa=1.74e-06 sb=5.97091e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=129030 $Y=53890 $D=28
M3547 3822 545 VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=1.02828e-13 pd=1.52e-06 ps=1.12945e-06 nrd=0.727273 nrs=0.531138 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=129470 $Y=54050 $D=28
M3548 3823 545 466 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=130430 $Y=54050 $D=28
M3549 466 545 3823 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=130910 $Y=54050 $D=28
M3550 3824 3822 466 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=131390 $Y=54050 $D=28
M3551 466 3822 3824 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-15 panw10=0 $X=131870 $Y=54050 $D=28
M3552 3825 17 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=11760 $Y=39490 $D=28
M3553 30 21 3825 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=12080 $Y=39490 $D=28
M3554 3826 21 30 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=12560 $Y=39490 $D=28
M3555 VSS 17 3826 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=12880 $Y=39490 $D=28
M3556 3827 17 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=13440 $Y=39490 $D=28
M3557 30 21 3827 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=13760 $Y=39490 $D=28
M3558 3828 14 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=12160 $Y=53890 $D=28
M3559 59 48 3828 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=12480 $Y=53890 $D=28
M3560 3829 48 59 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=12960 $Y=53890 $D=28
M3561 VSS 14 3829 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=13280 $Y=53890 $D=28
M3562 3830 14 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=13840 $Y=53890 $D=28
M3563 59 48 3830 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=14160 $Y=53890 $D=28
M3564 3831 34 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=14160 $Y=34190 $D=28
M3565 53 800 3831 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=14480 $Y=34190 $D=28
M3566 3832 800 53 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=14960 $Y=34090 $D=28
M3567 VSS 34 3832 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=15280 $Y=34090 $D=28
M3568 3833 34 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=15840 $Y=34090 $D=28
M3569 53 800 3833 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=16160 $Y=34090 $D=28
M3570 3834 73 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=26560 $Y=61090 $D=28
M3571 98 96 3834 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=26880 $Y=61090 $D=28
M3572 3835 96 98 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=27360 $Y=61090 $D=28
M3573 VSS 73 3835 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=27680 $Y=61090 $D=28
M3574 3836 73 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=28240 $Y=61090 $D=28
M3575 98 96 3836 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=28560 $Y=61090 $D=28
M3576 3837 148 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=38160 $Y=19790 $D=28
M3577 168 163 3837 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=38480 $Y=19790 $D=28
M3578 3838 163 168 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=38960 $Y=19690 $D=28
M3579 VSS 148 3838 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=39280 $Y=19690 $D=28
M3580 3839 148 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=39840 $Y=19690 $D=28
M3581 168 163 3839 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=40160 $Y=19690 $D=28
M3582 3840 148 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=42560 $Y=25090 $D=28
M3583 182 163 3840 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=42880 $Y=25090 $D=28
M3584 3841 163 182 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=43360 $Y=25090 $D=28
M3585 VSS 148 3841 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=43680 $Y=25090 $D=28
M3586 3842 148 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=44240 $Y=25090 $D=28
M3587 182 163 3842 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=44560 $Y=25090 $D=28
M3588 3843 143 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=47760 $Y=17890 $D=28
M3589 169 177 3843 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=48080 $Y=17890 $D=28
M3590 3844 177 169 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=48560 $Y=17890 $D=28
M3591 VSS 143 3844 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=48880 $Y=17890 $D=28
M3592 3845 143 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=49440 $Y=17890 $D=28
M3593 169 177 3845 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=49760 $Y=17890 $D=28
M3594 3846 278 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=64160 $Y=32290 $D=28
M3595 242 285 3846 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=64480 $Y=32290 $D=28
M3596 3847 285 242 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=64960 $Y=32290 $D=28
M3597 VSS 278 3847 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=65280 $Y=32290 $D=28
M3598 3848 278 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=65840 $Y=32290 $D=28
M3599 242 285 3848 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=66160 $Y=32290 $D=28
M3600 3849 213 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=64960 $Y=48590 $D=28
M3601 246 245 3849 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=65280 $Y=48590 $D=28
M3602 3850 245 246 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=65760 $Y=48490 $D=28
M3603 VSS 213 3850 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=66080 $Y=48490 $D=28
M3604 3851 213 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=66640 $Y=48490 $D=28
M3605 246 245 3851 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=66960 $Y=48490 $D=28
M3606 3852 278 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=72960 $Y=34190 $D=28
M3607 282 291 3852 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=73280 $Y=34190 $D=28
M3608 3853 291 282 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=73760 $Y=34090 $D=28
M3609 VSS 278 3853 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=74080 $Y=34090 $D=28
M3610 3854 278 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=74640 $Y=34090 $D=28
M3611 282 291 3854 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=74960 $Y=34090 $D=28
M3612 3855 308 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=78960 $Y=75490 $D=28
M3613 358 347 3855 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=79280 $Y=75490 $D=28
M3614 3856 347 358 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=79760 $Y=75490 $D=28
M3615 VSS 308 3856 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=80080 $Y=75490 $D=28
M3616 3857 308 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=80640 $Y=75490 $D=28
M3617 358 347 3857 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=80960 $Y=75490 $D=28
M3618 3858 301 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=79760 $Y=39490 $D=28
M3619 330 278 3858 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=80080 $Y=39490 $D=28
M3620 3859 278 330 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=80560 $Y=39490 $D=28
M3621 VSS 301 3859 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=80880 $Y=39490 $D=28
M3622 3860 301 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=81440 $Y=39490 $D=28
M3623 330 278 3860 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=81760 $Y=39490 $D=28
M3624 3861 392 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=105360 $Y=62990 $D=28
M3625 476 401 3861 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=105680 $Y=62990 $D=28
M3626 3862 401 476 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=106160 $Y=62890 $D=28
M3627 VSS 392 3862 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=106480 $Y=62890 $D=28
M3628 3863 392 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=107040 $Y=62890 $D=28
M3629 476 401 3863 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=107360 $Y=62890 $D=28
M3630 3864 427 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=114560 $Y=32290 $D=28
M3631 405 836 3864 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=114880 $Y=32290 $D=28
M3632 3865 836 405 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=115360 $Y=32290 $D=28
M3633 VSS 427 3865 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=115680 $Y=32290 $D=28
M3634 3866 427 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=116240 $Y=32290 $D=28
M3635 405 836 3866 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=116560 $Y=32290 $D=28
M3636 3867 490 VSS VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=2.304e-13 pd=9.2e-07 ps=2.08e-06 nrd=0.138889 nrs=0.444444 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=127360 $Y=75490 $D=28
M3637 496 473 3867 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3147e-13 as=7.2e-14 pd=1.10338e-06 ps=9.2e-07 nrd=0.253608 nrs=0.138889 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-15 panw10=0 $X=127680 $Y=75490 $D=28
M3638 3868 473 496 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.4973e-13 pd=1.02e-06 ps=1.25662e-06 nrd=0.121951 nrs=0.22268 sa=1.01024e-06 sb=1.52e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=128160 $Y=75490 $D=28
M3639 VSS 490 3868 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.98337e-13 as=8.2e-14 pd=1.39229e-06 ps=1.02e-06 nrd=0.29497 nrs=0.121951 sa=1.33024e-06 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=128480 $Y=75490 $D=28
M3640 3869 490 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.98337e-13 pd=1.02e-06 ps=1.39229e-06 nrd=0.121951 nrs=0.29497 sa=1.89024e-06 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=129040 $Y=75490 $D=28
M3641 496 473 3869 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=1.92927e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=129360 $Y=75490 $D=28
M3642 3870 216 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.6e-14 as=2.924e-13 pd=1.06e-06 ps=2.4e-06 nrd=0.116279 nrs=0.395349 sa=3.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=57230 $Y=41190 $D=28
M3643 284 206 3870 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=8.6e-14 pd=1.22e-06 ps=1.06e-06 nrd=0.209302 nrs=0.116279 sa=6.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=57550 $Y=41190 $D=28
M3644 3871 206 284 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.6e-14 as=1.548e-13 pd=1.06e-06 ps=1.22e-06 nrd=0.116279 nrs=0.209302 sa=1.14e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=58030 $Y=41190 $D=28
M3645 VSS 216 3871 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9522e-13 as=8.6e-14 pd=1.3502e-06 ps=1.06e-06 nrd=0.263953 nrs=0.116279 sa=1.46e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=58350 $Y=41190 $D=28
M3646 3872 216 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.6e-14 as=1.9522e-13 pd=1.06e-06 ps=1.3502e-06 nrd=0.116279 nrs=0.263953 sa=2e-06 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=58910 $Y=41190 $D=28
M3647 284 206 3872 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=8.6e-14 pd=1.22e-06 ps=1.06e-06 nrd=0.209302 nrs=0.116279 sa=2e-06 sb=1.33e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=59230 $Y=41190 $D=28
M3648 3873 206 284 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.6e-14 as=1.548e-13 pd=1.06e-06 ps=1.22e-06 nrd=0.116279 nrs=0.209302 sa=2e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=59710 $Y=41190 $D=28
M3649 VSS 216 3873 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.54411e-13 as=8.6e-14 pd=2.17263e-06 ps=1.06e-06 nrd=0.479192 nrs=0.116279 sa=2e-06 sb=5.3e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=60030 $Y=41190 $D=28
M3650 3874 278 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.6e-14 as=2.924e-13 pd=1.06e-06 ps=2.4e-06 nrd=0.116279 nrs=0.395349 sa=3.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=80030 $Y=33990 $D=28
M3651 232 304 3874 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=8.6e-14 pd=1.22e-06 ps=1.06e-06 nrd=0.209302 nrs=0.116279 sa=6.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=80350 $Y=33990 $D=28
M3652 3875 304 232 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.6e-14 as=1.548e-13 pd=1.06e-06 ps=1.22e-06 nrd=0.116279 nrs=0.209302 sa=1.14e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=80830 $Y=33990 $D=28
M3653 VSS 278 3875 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9522e-13 as=8.6e-14 pd=1.3502e-06 ps=1.06e-06 nrd=0.263953 nrs=0.116279 sa=1.46e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=81150 $Y=33990 $D=28
M3654 3876 278 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.6e-14 as=1.9522e-13 pd=1.06e-06 ps=1.3502e-06 nrd=0.116279 nrs=0.263953 sa=2e-06 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=81710 $Y=33990 $D=28
M3655 232 304 3876 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=8.6e-14 pd=1.22e-06 ps=1.06e-06 nrd=0.209302 nrs=0.116279 sa=2e-06 sb=1.33e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=82030 $Y=33990 $D=28
M3656 3877 304 232 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.6e-14 as=1.548e-13 pd=1.06e-06 ps=1.22e-06 nrd=0.116279 nrs=0.209302 sa=2e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=82510 $Y=33990 $D=28
M3657 VSS 278 3877 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.54411e-13 as=8.6e-14 pd=2.17263e-06 ps=1.06e-06 nrd=0.479192 nrs=0.116279 sa=2e-06 sb=5.3e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=82830 $Y=33990 $D=28
M3658 3878 460 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.6e-14 as=2.924e-13 pd=1.06e-06 ps=2.4e-06 nrd=0.116279 nrs=0.395349 sa=3.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=126430 $Y=62790 $D=28
M3659 846 443 3878 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=8.6e-14 pd=1.22e-06 ps=1.06e-06 nrd=0.209302 nrs=0.116279 sa=6.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=126750 $Y=62790 $D=28
M3660 3879 443 846 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.6e-14 as=1.548e-13 pd=1.06e-06 ps=1.22e-06 nrd=0.116279 nrs=0.209302 sa=1.14e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=127230 $Y=62790 $D=28
M3661 VSS 460 3879 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9522e-13 as=8.6e-14 pd=1.3502e-06 ps=1.06e-06 nrd=0.263953 nrs=0.116279 sa=1.46e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=127550 $Y=62790 $D=28
M3662 3880 460 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.6e-14 as=1.9522e-13 pd=1.06e-06 ps=1.3502e-06 nrd=0.116279 nrs=0.263953 sa=2e-06 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=128110 $Y=62790 $D=28
M3663 846 443 3880 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=8.6e-14 pd=1.22e-06 ps=1.06e-06 nrd=0.209302 nrs=0.116279 sa=2e-06 sb=1.33e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=128430 $Y=62790 $D=28
M3664 3881 443 846 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.6e-14 as=1.548e-13 pd=1.06e-06 ps=1.22e-06 nrd=0.116279 nrs=0.209302 sa=2e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=128910 $Y=62790 $D=28
M3665 VSS 460 3881 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.54411e-13 as=8.6e-14 pd=2.17263e-06 ps=1.06e-06 nrd=0.479192 nrs=0.116279 sa=2e-06 sb=5.3e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=129230 $Y=62790 $D=28
M3666 VSS 228 3882 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.5538e-13 as=2.752e-13 pd=1.23685e-06 ps=2.36e-06 nrd=0.210086 nrs=0.372093 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=56840 $Y=55590 $D=28
M3667 211 218 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.6622e-13 pd=1.28e-06 ps=1.32315e-06 nrd=0.195652 nrs=0.196385 sa=7.6087e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=57320 $Y=55590 $D=28
M3668 VSS 3882 211 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.24087e-06 sb=1.72e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=57800 $Y=55590 $D=28
M3669 211 3882 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.72087e-06 sb=1.24e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=58280 $Y=55590 $D=28
M3670 VSS 218 211 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.15112e-13 as=1.656e-13 pd=1.97143e-06 ps=1.28e-06 nrd=0.490444 nrs=0.195652 sa=1.97652e-06 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=58760 $Y=55590 $D=28
M3671 VSS 466 3886 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.5538e-13 as=2.752e-13 pd=1.23685e-06 ps=2.36e-06 nrd=0.210086 nrs=0.372093 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=124040 $Y=53950 $D=28
M3672 475 485 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.6622e-13 pd=1.28e-06 ps=1.32315e-06 nrd=0.195652 nrs=0.196385 sa=7.6087e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=124520 $Y=53890 $D=28
M3673 VSS 3886 475 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.24087e-06 sb=1.72e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=125000 $Y=53890 $D=28
M3674 475 3886 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.72087e-06 sb=1.24e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=125480 $Y=53890 $D=28
M3675 VSS 485 475 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.15112e-13 as=1.656e-13 pd=1.97143e-06 ps=1.28e-06 nrd=0.490444 nrs=0.195652 sa=1.97652e-06 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=125960 $Y=53890 $D=28
M3676 3890 8 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=2.112e-13 pd=1.02e-06 ps=1.96e-06 nrd=0.272727 nrs=0.484848 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=9000 $Y=39490 $D=28
M3677 VSS 17 3890 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.77135e-13 as=1.188e-13 pd=1.19935e-06 ps=1.02e-06 nrd=0.406647 nrs=0.272727 sa=8e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=9480 $Y=39490 $D=28
M3678 14 3890 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.46916e-13 pd=1.28e-06 ps=1.67183e-06 nrd=0.195652 nrs=0.291725 sa=1.12043e-06 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=10100 $Y=39490 $D=28
M3679 VSS 3890 14 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=1.60043e-06 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=10580 $Y=39490 $D=28
M3680 3892 156 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=2.112e-13 pd=1.02e-06 ps=1.96e-06 nrd=0.272727 nrs=0.484848 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=36600 $Y=53890 $D=28
M3681 VSS 146 3892 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.77135e-13 as=1.188e-13 pd=1.19935e-06 ps=1.02e-06 nrd=0.406647 nrs=0.272727 sa=8e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=37080 $Y=53890 $D=28
M3682 138 3892 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.46916e-13 pd=1.28e-06 ps=1.67183e-06 nrd=0.195652 nrs=0.291725 sa=1.12043e-06 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=37700 $Y=53890 $D=28
M3683 VSS 3892 138 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=1.60043e-06 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=38180 $Y=53890 $D=28
M3684 3894 146 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=2.112e-13 pd=1.02e-06 ps=1.96e-06 nrd=0.272727 nrs=0.484848 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=39800 $Y=55850 $D=28
M3685 VSS 156 3894 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.77135e-13 as=1.188e-13 pd=1.19935e-06 ps=1.02e-06 nrd=0.406647 nrs=0.272727 sa=8e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=40280 $Y=55850 $D=28
M3686 160 3894 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.46916e-13 pd=1.28e-06 ps=1.67183e-06 nrd=0.195652 nrs=0.291725 sa=1.12043e-06 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=40900 $Y=55590 $D=28
M3687 VSS 3894 160 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=1.60043e-06 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=41380 $Y=55590 $D=28
M3688 3896 248 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=2.112e-13 pd=1.02e-06 ps=1.96e-06 nrd=0.272727 nrs=0.484848 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=75800 $Y=55850 $D=28
M3689 VSS 239 3896 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.77135e-13 as=1.188e-13 pd=1.19935e-06 ps=1.02e-06 nrd=0.406647 nrs=0.272727 sa=8e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=76280 $Y=55850 $D=28
M3690 315 3896 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.46916e-13 pd=1.28e-06 ps=1.67183e-06 nrd=0.195652 nrs=0.291725 sa=1.12043e-06 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=76900 $Y=55590 $D=28
M3691 VSS 3896 315 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=1.60043e-06 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=77380 $Y=55590 $D=28
M3692 3898 463 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=2.112e-13 pd=1.02e-06 ps=1.96e-06 nrd=0.272727 nrs=0.484848 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=121400 $Y=53890 $D=28
M3693 VSS 457 3898 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.77135e-13 as=1.188e-13 pd=1.19935e-06 ps=1.02e-06 nrd=0.406647 nrs=0.272727 sa=8e-07 sb=1.44e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=121880 $Y=53890 $D=28
M3694 460 3898 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.46916e-13 pd=1.28e-06 ps=1.67183e-06 nrd=0.195652 nrs=0.291725 sa=1.12043e-06 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=122500 $Y=53890 $D=28
M3695 VSS 3898 460 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=1.60043e-06 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=122980 $Y=53890 $D=28
M3696 799 40 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=2.112e-13 pd=1.02e-06 ps=1.96e-06 nrd=0.272727 nrs=0.484848 sa=3.2e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=14090 $Y=19850 $D=28
M3697 VSS 40 799 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.772e-13 as=1.188e-13 pd=2.16e-06 ps=1.02e-06 nrd=0.636364 nrs=0.272727 sa=8e-07 sb=4.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=14570 $Y=19850 $D=28
M3698 177 188 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=2.112e-13 pd=1.02e-06 ps=1.96e-06 nrd=0.272727 nrs=0.484848 sa=3.2e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=46090 $Y=17890 $D=28
M3699 VSS 188 177 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.772e-13 as=1.188e-13 pd=2.16e-06 ps=1.02e-06 nrd=0.636364 nrs=0.272727 sa=8e-07 sb=4.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=46570 $Y=17890 $D=28
M3700 377 368 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=2.112e-13 pd=1.02e-06 ps=1.96e-06 nrd=0.272727 nrs=0.484848 sa=3.2e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=94490 $Y=17890 $D=28
M3701 VSS 368 377 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.772e-13 as=1.188e-13 pd=2.16e-06 ps=1.02e-06 nrd=0.636364 nrs=0.272727 sa=8e-07 sb=4.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=94970 $Y=17890 $D=28
M3702 836 441 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=2.112e-13 pd=1.02e-06 ps=1.96e-06 nrd=0.272727 nrs=0.484848 sa=3.2e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=112890 $Y=32290 $D=28
M3703 VSS 441 836 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.772e-13 as=1.188e-13 pd=2.16e-06 ps=1.02e-06 nrd=0.636364 nrs=0.272727 sa=8e-07 sb=4.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=113370 $Y=32290 $D=28
M3704 467 432 VSS VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=2.112e-13 pd=1.02e-06 ps=1.96e-06 nrd=0.272727 nrs=0.484848 sa=3.2e-07 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=119290 $Y=61090 $D=28
M3705 VSS 432 467 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.772e-13 as=1.188e-13 pd=2.16e-06 ps=1.02e-06 nrd=0.636364 nrs=0.272727 sa=8e-07 sb=4.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=119770 $Y=61090 $D=28
M3706 VSS 910 3902 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.72e-13 as=2.944e-13 pd=1.63e-06 ps=2.48e-06 nrd=0.203214 nrs=0.347826 sa=3.2e-07 sb=1.17739e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=110410 $Y=46690 $D=28
M3707 3900 3902 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16285e-13 as=1.19652e-13 pd=1.08475e-06 ps=1.13391e-06 nrd=0.283898 nrs=0.29212 sa=7.6e-07 sb=1.38125e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=110850 $Y=46690 $D=28
M3708 3904 3901 3900 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62491e-13 as=9.81153e-14 pd=1.30091e-06 ps=9.15254e-07 nrd=0.557239 nrs=0.336472 sa=1.24e-06 sb=1.42222e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=111330 $Y=46690 $D=28
M3709 3901 3900 3904 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.00696e-14 as=1.02309e-13 pd=6.94783e-07 ps=8.19091e-07 nrd=0.606138 nrs=0.885027 sa=1.88e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=111970 $Y=46690 $D=28
M3710 VSS 436 3901 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.61391e-13 as=1.1953e-13 pd=1.72739e-06 ps=1.18522e-06 nrd=0.47976 nrs=0.355322 sa=1.28828e-06 sb=1.26086e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=9.6e-15 panw9=0 panw10=0 $X=112450 $Y=46690 $D=28
M3711 3901 436 VSS VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.8e-14 as=9.46087e-14 pd=7.4e-07 ps=1.01261e-06 nrd=0.588235 nrs=0.818414 sa=2e-06 sb=1.89088e-06 sd=0 panw1=0 panw2=3.5e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.3e-15 panw8=0 panw9=0 panw10=0 $X=112890 $Y=46690 $D=28
M3712 3906 3902 3901 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.89273e-14 as=6.8e-14 pd=6.95455e-07 ps=7.4e-07 nrd=0.596257 nrs=0.588235 sa=2e-06 sb=1.75206e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=113410 $Y=46690 $D=28
M3713 3902 3901 3906 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.89377e-13 as=1.09473e-13 pd=1.44419e-06 ps=1.10455e-06 nrd=0.64944 nrs=0.375421 sa=1.36296e-06 sb=9.75e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=113890 $Y=46690 $D=28
M3714 3905 3906 3902 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.76e-14 as=1.12223e-13 pd=6.8e-07 ps=8.55814e-07 nrd=0.5625 nrs=1.09593 sa=1.76094e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=114570 $Y=46640 $D=28
M3715 3903 3904 3905 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.42e-13 as=5.76e-14 pd=1.37e-06 ps=6.8e-07 nrd=1.38672 nrs=0.5625 sa=1.83594e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=115050 $Y=46640 $D=28
M3716 VSS 451 3903 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.0176e-13 as=1.42e-13 pd=1.01333e-06 ps=1.37e-06 nrd=0.99375 nrs=1.38672 sa=3.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=6e-15 panw9=3.24e-14 panw10=0 $X=115570 $Y=47290 $D=28
M3717 3907 451 3904 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.12e-14 as=1.088e-13 pd=7e-07 ps=1.32e-06 nrd=0.529412 nrs=0.941176 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.32e-14 panw8=0 panw9=0 panw10=0 $X=116290 $Y=46760 $D=28
M3718 3906 3903 3907 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=6.12e-14 pd=1.32e-06 ps=7e-07 nrd=0.941176 nrs=0.529412 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.32e-14 panw8=0 panw9=0 panw10=0 $X=116770 $Y=46760 $D=28
M3719 VSS 3905 480 VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.584e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.366213 sa=3.07619e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=117690 $Y=46760 $D=28
M3720 457 3907 VSS VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=7.87619e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=118170 $Y=46760 $D=28
M3721 VSS 839 3910 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.72e-13 as=2.944e-13 pd=1.63e-06 ps=2.48e-06 nrd=0.203214 nrs=0.347826 sa=3.2e-07 sb=1.17739e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=118410 $Y=41190 $D=28
M3722 3908 3910 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16285e-13 as=1.19652e-13 pd=1.08475e-06 ps=1.13391e-06 nrd=0.283898 nrs=0.29212 sa=7.6e-07 sb=1.38125e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=118850 $Y=41470 $D=28
M3723 3912 3909 3908 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62491e-13 as=9.81153e-14 pd=1.30091e-06 ps=9.15254e-07 nrd=0.557239 nrs=0.336472 sa=1.24e-06 sb=1.42222e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=119330 $Y=41570 $D=28
M3724 3909 3908 3912 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.00696e-14 as=1.02309e-13 pd=6.94783e-07 ps=8.19091e-07 nrd=0.606138 nrs=0.885027 sa=1.88e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=119970 $Y=41770 $D=28
M3725 VSS 444 3909 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.61391e-13 as=1.1953e-13 pd=1.72739e-06 ps=1.18522e-06 nrd=0.47976 nrs=0.355322 sa=1.28828e-06 sb=1.26086e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=9.6e-15 panw9=0 panw10=0 $X=120450 $Y=41530 $D=28
M3726 3909 444 VSS VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.8e-14 as=9.46087e-14 pd=7.4e-07 ps=1.01261e-06 nrd=0.588235 nrs=0.818414 sa=2e-06 sb=1.89088e-06 sd=0 panw1=0 panw2=3.5e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.3e-15 panw8=0 panw9=0 panw10=0 $X=120890 $Y=41770 $D=28
M3727 3914 3910 3909 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.89273e-14 as=6.8e-14 pd=6.95455e-07 ps=7.4e-07 nrd=0.596257 nrs=0.588235 sa=2e-06 sb=1.75206e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=121410 $Y=41770 $D=28
M3728 3910 3909 3914 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.89377e-13 as=1.09473e-13 pd=1.44419e-06 ps=1.10455e-06 nrd=0.64944 nrs=0.375421 sa=1.36296e-06 sb=9.75e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=121890 $Y=41570 $D=28
M3729 3913 3914 3910 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.76e-14 as=1.12223e-13 pd=6.8e-07 ps=8.55814e-07 nrd=0.5625 nrs=1.09593 sa=1.76094e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=122570 $Y=41840 $D=28
M3730 3911 3912 3913 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.42e-13 as=5.76e-14 pd=1.37e-06 ps=6.8e-07 nrd=1.38672 nrs=0.5625 sa=1.83594e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=123050 $Y=41840 $D=28
M3731 VSS 403 3911 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.0176e-13 as=1.42e-13 pd=1.01333e-06 ps=1.37e-06 nrd=0.99375 nrs=1.38672 sa=3.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=6e-15 panw9=3.24e-14 panw10=1.2e-14 $X=123570 $Y=41190 $D=28
M3732 3915 403 3912 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.12e-14 as=1.088e-13 pd=7e-07 ps=1.32e-06 nrd=0.529412 nrs=0.941176 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.32e-14 panw8=0 panw9=0 panw10=0 $X=124290 $Y=41700 $D=28
M3733 3914 3911 3915 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=6.12e-14 pd=1.32e-06 ps=7e-07 nrd=0.941176 nrs=0.529412 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.32e-14 panw8=0 panw9=0 panw10=0 $X=124770 $Y=41700 $D=28
M3734 VSS 3913 470 VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.584e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.366213 sa=3.07619e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=125690 $Y=41200 $D=28
M3735 845 3915 VSS VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=7.87619e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=126170 $Y=41200 $D=28
M3736 VSS 189 3916 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.952e-13 pd=9.7e-07 ps=1.86e-06 nrd=0.295082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=40040 $Y=61090 $D=28
M3737 3916 174 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=40520 $Y=61090 $D=28
M3738 VSS 174 3916 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30296e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.350164 nrs=0.295082 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=41000 $Y=61090 $D=28
M3739 3916 189 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.30296e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.350164 sa=1.72e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=41440 $Y=61090 $D=28
M3740 152 180 3916 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=41920 $Y=61090 $D=28
M3741 3916 151 152 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=42400 $Y=61090 $D=28
M3742 152 151 3916 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=42880 $Y=61090 $D=28
M3743 3916 180 152 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=43360 $Y=61090 $D=28
M3744 VSS 203 3921 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.952e-13 pd=9.7e-07 ps=1.86e-06 nrd=0.295082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=41240 $Y=19900 $D=28
M3745 3921 182 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=41720 $Y=19900 $D=28
M3746 VSS 182 3921 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30296e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.350164 nrs=0.295082 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=42200 $Y=19900 $D=28
M3747 3921 203 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.30296e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.350164 sa=1.72e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=42640 $Y=19900 $D=28
M3748 173 148 3921 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=43120 $Y=19900 $D=28
M3749 3921 165 173 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=43600 $Y=19900 $D=28
M3750 173 165 3921 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=44080 $Y=19900 $D=28
M3751 3921 148 173 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=44560 $Y=19900 $D=28
M3752 VSS 179 3926 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.952e-13 pd=9.7e-07 ps=1.86e-06 nrd=0.295082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=43640 $Y=63100 $D=28
M3753 3926 189 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=44120 $Y=63100 $D=28
M3754 VSS 189 3926 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30296e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.350164 nrs=0.295082 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=44600 $Y=63100 $D=28
M3755 3926 179 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.30296e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.350164 sa=1.72e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=45040 $Y=63100 $D=28
M3756 894 174 3926 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=45520 $Y=63100 $D=28
M3757 3926 151 894 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=46000 $Y=63100 $D=28
M3758 894 151 3926 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=46480 $Y=63100 $D=28
M3759 3926 174 894 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=46960 $Y=63100 $D=28
M3760 VSS 148 3931 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.952e-13 pd=9.7e-07 ps=1.86e-06 nrd=0.295082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=45240 $Y=41500 $D=28
M3761 3931 185 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=45720 $Y=41500 $D=28
M3762 VSS 185 3931 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30296e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.350164 nrs=0.295082 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=46200 $Y=41500 $D=28
M3763 3931 148 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.30296e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.350164 sa=1.72e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=46640 $Y=41500 $D=28
M3764 812 166 3931 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=47120 $Y=41500 $D=28
M3765 3931 168 812 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=47600 $Y=41500 $D=28
M3766 812 168 3931 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=48080 $Y=41500 $D=28
M3767 3931 166 812 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=48560 $Y=41500 $D=28
M3768 VSS 148 3936 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.952e-13 pd=9.7e-07 ps=1.86e-06 nrd=0.295082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=50840 $Y=53890 $D=28
M3769 3936 200 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=51320 $Y=53890 $D=28
M3770 VSS 200 3936 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30296e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.350164 nrs=0.295082 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=51800 $Y=53890 $D=28
M3771 3936 148 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.30296e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.350164 sa=1.72e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=52240 $Y=53890 $D=28
M3772 210 185 3936 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=52720 $Y=53890 $D=28
M3773 3936 168 210 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=53200 $Y=53890 $D=28
M3774 210 168 3936 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=53680 $Y=53890 $D=28
M3775 3936 185 210 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=54160 $Y=53890 $D=28
M3776 VSS 203 3941 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.952e-13 pd=9.7e-07 ps=1.86e-06 nrd=0.295082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=54840 $Y=27100 $D=28
M3777 3941 148 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=55320 $Y=27100 $D=28
M3778 VSS 148 3941 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30296e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.350164 nrs=0.295082 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=55800 $Y=27100 $D=28
M3779 3941 203 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.30296e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.350164 sa=1.72e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=56240 $Y=27100 $D=28
M3780 227 217 3941 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=56720 $Y=27100 $D=28
M3781 3941 198 227 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=57200 $Y=27100 $D=28
M3782 227 198 3941 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=57680 $Y=27100 $D=28
M3783 3941 217 227 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=58160 $Y=27100 $D=28
M3784 VSS 291 3946 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.952e-13 pd=9.7e-07 ps=1.86e-06 nrd=0.295082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=67240 $Y=41500 $D=28
M3785 3946 820 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=67720 $Y=41500 $D=28
M3786 VSS 820 3946 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30296e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.350164 nrs=0.295082 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=68200 $Y=41500 $D=28
M3787 3946 291 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.30296e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.350164 sa=1.72e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=68640 $Y=41500 $D=28
M3788 215 267 3946 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=69120 $Y=41500 $D=28
M3789 3946 232 215 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=69600 $Y=41500 $D=28
M3790 215 232 3946 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=70080 $Y=41500 $D=28
M3791 3946 267 215 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=70560 $Y=41500 $D=28
M3792 VSS 213 3951 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.952e-13 pd=9.7e-07 ps=1.86e-06 nrd=0.295082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=68840 $Y=55900 $D=28
M3793 3951 280 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=69320 $Y=55900 $D=28
M3794 VSS 280 3951 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30296e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.350164 nrs=0.295082 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=69800 $Y=55900 $D=28
M3795 3951 213 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.30296e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.350164 sa=1.72e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=70240 $Y=55900 $D=28
M3796 266 246 3951 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=70720 $Y=55900 $D=28
M3797 3951 255 266 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=71200 $Y=55900 $D=28
M3798 266 255 3951 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=71680 $Y=55900 $D=28
M3799 3951 246 266 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=72160 $Y=55900 $D=28
M3800 VSS 319 3956 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.952e-13 pd=9.7e-07 ps=1.86e-06 nrd=0.295082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=87240 $Y=41500 $D=28
M3801 3956 336 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=87720 $Y=41500 $D=28
M3802 VSS 336 3956 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30296e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.350164 nrs=0.295082 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=88200 $Y=41500 $D=28
M3803 3956 319 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.30296e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.350164 sa=1.72e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=88640 $Y=41500 $D=28
M3804 320 313 3956 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=89120 $Y=41500 $D=28
M3805 3956 330 320 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=89600 $Y=41500 $D=28
M3806 320 330 3956 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=90080 $Y=41500 $D=28
M3807 3956 313 320 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=90560 $Y=41500 $D=28
M3808 VSS 419 3961 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.952e-13 pd=9.7e-07 ps=1.86e-06 nrd=0.295082 nrs=0.52459 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=114040 $Y=41500 $D=28
M3809 3961 410 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=114520 $Y=41500 $D=28
M3810 VSS 410 3961 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30296e-13 as=1.098e-13 pd=1.32573e-06 ps=9.7e-07 nrd=0.350164 nrs=0.295082 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=115000 $Y=41500 $D=28
M3811 3961 419 VSS VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.30296e-13 pd=9.7e-07 ps=1.32573e-06 nrd=0.295082 nrs=0.350164 sa=1.72e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=115440 $Y=41500 $D=28
M3812 446 400 3961 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=115920 $Y=41500 $D=28
M3813 3961 416 446 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=116400 $Y=41500 $D=28
M3814 446 416 3961 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.098e-13 as=1.098e-13 pd=9.7e-07 ps=9.7e-07 nrd=0.295082 nrs=0.295082 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=116880 $Y=41500 $D=28
M3815 3961 400 446 VSS lpnfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.952e-13 as=1.098e-13 pd=1.86e-06 ps=9.7e-07 nrd=0.52459 nrs=0.295082 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=117360 $Y=41500 $D=28
M3816 3973 3966 3967 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96060 $Y=46710 $D=28
M3817 3975 357 3973 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96380 $Y=46710 $D=28
M3818 VSS 329 3975 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=96700 $Y=46710 $D=28
M3819 VSS clk 3966 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=97680 $Y=46860 $D=28
M3820 3969 3966 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=98190 $Y=46860 $D=28
M3821 3977 3969 3967 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=99210 $Y=46790 $D=28
M3822 3978 3968 3977 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=99530 $Y=46790 $D=28
M3823 VSS 329 3978 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=99850 $Y=46790 $D=28
M3824 3968 3967 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=100310 $Y=46930 $D=28
M3825 3970 3969 3968 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=100870 $Y=46930 $D=28
M3826 3980 3966 3970 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=101430 $Y=46690 $D=28
M3827 VSS 3972 3980 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.27475e-14 as=2e-14 pd=5.0303e-07 ps=4e-07 nrd=1.81869 nrs=0.5 sa=6.6e-07 sb=1.08e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=101750 $Y=46690 $D=28
M3828 3981 329 VSS VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.2e-14 as=1.16396e-13 pd=5.2e-07 ps=8.04848e-07 nrd=0.3125 nrs=1.13668 sa=7.775e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=102190 $Y=46690 $D=28
M3829 3972 3970 3981 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.024e-13 as=3.2e-14 pd=1.28e-06 ps=5.2e-07 nrd=1 nrs=0.3125 sa=1.0975e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=102510 $Y=46690 $D=28
M3830 3971 3972 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.27475e-14 pd=1.28e-06 ps=5.0303e-07 nrd=2.36 nrs=1.81869 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=102830 $Y=47410 $D=28
M3831 VSS 3971 942 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.32327e-13 as=1.472e-13 pd=1.24967e-06 ps=1.56e-06 nrd=0.625362 nrs=0.695652 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=103790 $Y=46690 $D=28
M3832 359 3972 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.32327e-13 pd=1.56e-06 ps=1.24967e-06 nrd=0.695652 nrs=0.625362 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=104270 $Y=46690 $D=28
M3833 3989 3982 3983 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=103260 $Y=56290 $D=28
M3834 3991 369 3989 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=103580 $Y=56290 $D=28
M3835 VSS 374 3991 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=103900 $Y=56290 $D=28
M3836 VSS clk 3982 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=104880 $Y=56040 $D=28
M3837 3985 3982 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=105390 $Y=56140 $D=28
M3838 3993 3985 3983 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=106410 $Y=56210 $D=28
M3839 3994 3984 3993 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=106730 $Y=56210 $D=28
M3840 VSS 374 3994 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=107050 $Y=56210 $D=28
M3841 3984 3983 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=107510 $Y=56070 $D=28
M3842 3986 3985 3984 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=108070 $Y=56070 $D=28
M3843 3996 3982 3986 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=108630 $Y=56310 $D=28
M3844 VSS 3988 3996 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.27475e-14 as=2e-14 pd=5.0303e-07 ps=4e-07 nrd=1.81869 nrs=0.5 sa=6.6e-07 sb=1.08e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=108950 $Y=56310 $D=28
M3845 3997 374 VSS VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.2e-14 as=1.16396e-13 pd=5.2e-07 ps=8.04848e-07 nrd=0.3125 nrs=1.13668 sa=7.775e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=109390 $Y=56190 $D=28
M3846 3988 3986 3997 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.024e-13 as=3.2e-14 pd=1.28e-06 ps=5.2e-07 nrd=1 nrs=0.3125 sa=1.0975e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=109710 $Y=56190 $D=28
M3847 3987 3988 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.27475e-14 pd=1.28e-06 ps=5.0303e-07 nrd=2.36 nrs=1.81869 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=110030 $Y=55590 $D=28
M3848 VSS 3987 837 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.32327e-13 as=1.472e-13 pd=1.24967e-06 ps=1.56e-06 nrd=0.625362 nrs=0.695652 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=110990 $Y=56050 $D=28
M3849 418 3988 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.32327e-13 pd=1.56e-06 ps=1.24967e-06 nrd=0.695652 nrs=0.625362 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=111470 $Y=56050 $D=28
M3850 4005 3998 3999 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=112060 $Y=53910 $D=28
M3851 4007 835 4005 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=112380 $Y=53910 $D=28
M3852 VSS 425 4007 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=112700 $Y=53910 $D=28
M3853 VSS clk 3998 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=113680 $Y=54060 $D=28
M3854 4001 3998 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.56667e-14 pd=1.28e-06 ps=7.48718e-07 nrd=2.36 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=114190 $Y=54060 $D=28
M3855 4009 4001 3999 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.23e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=115210 $Y=53990 $D=28
M3856 4010 4000 4009 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=9.16e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=115530 $Y=53990 $D=28
M3857 VSS 425 4010 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.132e-13 as=2e-14 pd=1.32e-06 ps=4e-07 nrd=2.83 nrs=0.5 sa=1e-06 sb=5.96e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=115850 $Y=53990 $D=28
M3858 4000 3999 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.52e-14 as=1.132e-13 pd=7.2e-07 ps=1.32e-06 nrd=1.38 nrs=2.83 sa=6.2e-07 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=116310 $Y=54130 $D=28
M3859 4002 4001 4000 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=5.52e-14 pd=9.6e-07 ps=7.2e-07 nrd=2.16 nrs=1.38 sa=1.174e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=116870 $Y=54130 $D=28
M3860 4012 3998 4002 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=8.64e-14 pd=4e-07 ps=9.6e-07 nrd=0.5 nrs=2.16 sa=3.4e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=117430 $Y=53890 $D=28
M3861 VSS 4004 4012 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.27475e-14 as=2e-14 pd=5.0303e-07 ps=4e-07 nrd=1.81869 nrs=0.5 sa=6.6e-07 sb=1.08e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=117750 $Y=53890 $D=28
M3862 4013 425 VSS VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.2e-14 as=1.16396e-13 pd=5.2e-07 ps=8.04848e-07 nrd=0.3125 nrs=1.13668 sa=7.775e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=118190 $Y=53890 $D=28
M3863 4004 4002 4013 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.024e-13 as=3.2e-14 pd=1.28e-06 ps=5.2e-07 nrd=1 nrs=0.3125 sa=1.0975e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=118510 $Y=53890 $D=28
M3864 4003 4004 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.44e-14 as=7.27475e-14 pd=1.28e-06 ps=5.0303e-07 nrd=2.36 nrs=1.81869 sa=1.14e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.4e-14 panw10=0 $X=118830 $Y=54610 $D=28
M3865 VSS 4003 943 VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.32327e-13 as=1.472e-13 pd=1.24967e-06 ps=1.56e-06 nrd=0.625362 nrs=0.695652 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=119790 $Y=53890 $D=28
M3866 452 4004 VSS VSS lpnfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.472e-13 as=1.32327e-13 pd=1.56e-06 ps=1.24967e-06 nrd=0.695652 nrs=0.625362 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=120270 $Y=53890 $D=28
M3867 4015 93 VSS VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.062e-13 as=1.888e-13 pd=9.5e-07 ps=1.82e-06 nrd=0.305085 nrs=0.542373 sa=3.2e-07 sb=1.14305e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=8810 $Y=25250 $D=28
M3868 VSS 93 4015 VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22021e-13 as=1.062e-13 pd=1.28489e-06 ps=9.5e-07 nrd=0.350534 nrs=0.305085 sa=8e-07 sb=6.63051e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=9290 $Y=25250 $D=28
M3869 4014 93 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=9.92711e-14 pd=1.6e-06 ps=1.04533e-06 nrd=0.666667 nrs=0.430864 sa=1.24e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=9730 $Y=25250 $D=28
M3870 VSS 4014 4016 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47609e-13 as=1.696e-13 pd=1.16284e-06 ps=1.7e-06 nrd=0.525486 nrs=0.603774 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=10770 $Y=25250 $D=28
M3871 4016 4014 VSS VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.54e-14 as=1.47609e-13 pd=8.9e-07 ps=1.16284e-06 nrd=0.339623 nrs=0.525486 sa=8.8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=11330 $Y=25250 $D=28
M3872 4017 90 4016 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.34138e-13 as=9.54e-14 pd=1.07927e-06 ps=8.9e-07 nrd=0.47753 nrs=0.339623 sa=1.36e-06 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=11810 $Y=25250 $D=28
M3873 4016 90 4017 VSS lpnfet w=5.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.824e-13 as=1.44262e-13 pd=1.78e-06 ps=1.16073e-06 nrd=0.561404 nrs=0.444019 sa=1.81053e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=12370 $Y=25210 $D=28
M3874 4017 4018 4015 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=13310 $Y=25140 $D=28
M3875 4015 4018 4017 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=13790 $Y=25140 $D=28
M3876 4020 90 4015 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=14270 $Y=25140 $D=28
M3877 4015 90 4020 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=14750 $Y=25140 $D=28
M3878 4016 4018 4020 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21e-13 as=3.016e-13 pd=9.9e-07 ps=2.56e-06 nrd=0.4 nrs=0.997025 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=15790 $Y=25090 $D=28
M3879 4020 4018 4016 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.016e-13 as=1.21e-13 pd=2.56e-06 ps=9.9e-07 nrd=0.997025 nrs=0.4 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=16350 $Y=25090 $D=28
M3880 VSS 90 4018 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.18002e-13 as=3.464e-13 pd=1.3493e-06 ps=2.52e-06 nrd=0.377428 nrs=0.599723 sa=4.3e-07 sb=1.71605e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=17540 $Y=25160 $D=28
M3881 4018 90 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45741e-13 as=2.18002e-13 pd=1.25176e-06 ps=1.3493e-06 nrd=0.252322 nrs=0.377428 sa=1.09e-06 sb=1.51632e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=18200 $Y=25160 $D=28
M3882 4019 4017 4018 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.235e-13 as=1.15059e-13 pd=1.07e-06 ps=9.88235e-07 nrd=0.343056 nrs=0.319608 sa=1.57e-06 sb=1.79e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=18680 $Y=25160 $D=28
M3883 4022 4020 4019 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.235e-13 pd=9.6e-07 ps=1.07e-06 nrd=0.3 nrs=0.343056 sa=1.80167e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=19200 $Y=25090 $D=28
M3884 4023 4017 4022 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.85767e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=19680 $Y=25090 $D=28
M3885 4021 4020 4023 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10571e-13 as=1.08e-13 pd=9.71429e-07 ps=9.6e-07 nrd=0.307143 nrs=0.3 sa=1.91367e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=20160 $Y=25090 $D=28
M3886 VSS 4022 4021 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.63084e-13 as=1.21629e-13 pd=1.15677e-06 ps=1.06857e-06 nrd=0.374389 nrs=0.279221 sa=1.81515e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=20640 $Y=25090 $D=28
M3887 4022 66 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.27329e-13 pd=2.48e-06 ps=1.61247e-06 nrd=0.347826 nrs=0.268583 sa=1.46022e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=21200 $Y=25090 $D=28
M3888 VSS 4019 17 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=22160 $Y=25090 $D=28
M3889 39 4023 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=22640 $Y=25090 $D=28
M3890 4025 150 VSS VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.062e-13 as=1.888e-13 pd=9.5e-07 ps=1.82e-06 nrd=0.305085 nrs=0.542373 sa=3.2e-07 sb=1.14305e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=8810 $Y=41360 $D=28
M3891 VSS 150 4025 VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22021e-13 as=1.062e-13 pd=1.28489e-06 ps=9.5e-07 nrd=0.350534 nrs=0.305085 sa=8e-07 sb=6.63051e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=9290 $Y=41360 $D=28
M3892 4024 150 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=9.92711e-14 pd=1.6e-06 ps=1.04533e-06 nrd=0.666667 nrs=0.430864 sa=1.24e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=9730 $Y=41470 $D=28
M3893 VSS 4024 4026 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47609e-13 as=1.696e-13 pd=1.16284e-06 ps=1.7e-06 nrd=0.525486 nrs=0.603774 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=10770 $Y=41420 $D=28
M3894 4026 4024 VSS VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.54e-14 as=1.47609e-13 pd=8.9e-07 ps=1.16284e-06 nrd=0.339623 nrs=0.525486 sa=8.8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=11330 $Y=41420 $D=28
M3895 4027 53 4026 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.34138e-13 as=9.54e-14 pd=1.07927e-06 ps=8.9e-07 nrd=0.47753 nrs=0.339623 sa=1.36e-06 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=11810 $Y=41420 $D=28
M3896 4026 53 4027 VSS lpnfet w=5.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.824e-13 as=1.44262e-13 pd=1.78e-06 ps=1.16073e-06 nrd=0.561404 nrs=0.444019 sa=1.81053e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=12370 $Y=41420 $D=28
M3897 4027 4028 4025 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=13310 $Y=41510 $D=28
M3898 4025 4028 4027 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=13790 $Y=41510 $D=28
M3899 4030 53 4025 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=14270 $Y=41510 $D=28
M3900 4025 53 4030 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=14750 $Y=41510 $D=28
M3901 4026 4028 4030 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21e-13 as=3.016e-13 pd=9.9e-07 ps=2.56e-06 nrd=0.4 nrs=0.997025 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=15790 $Y=41560 $D=28
M3902 4030 4028 4026 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.016e-13 as=1.21e-13 pd=2.56e-06 ps=9.9e-07 nrd=0.997025 nrs=0.4 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=16350 $Y=41560 $D=28
M3903 VSS 53 4028 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.18002e-13 as=3.464e-13 pd=1.3493e-06 ps=2.52e-06 nrd=0.377428 nrs=0.599723 sa=4.3e-07 sb=1.71605e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=17540 $Y=41280 $D=28
M3904 4028 53 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45741e-13 as=2.18002e-13 pd=1.25176e-06 ps=1.3493e-06 nrd=0.252322 nrs=0.377428 sa=1.09e-06 sb=1.51632e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=18200 $Y=41280 $D=28
M3905 4029 4027 4028 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.235e-13 as=1.15059e-13 pd=1.07e-06 ps=9.88235e-07 nrd=0.343056 nrs=0.319608 sa=1.57e-06 sb=1.79e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=18680 $Y=41440 $D=28
M3906 4032 4030 4029 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.235e-13 pd=9.6e-07 ps=1.07e-06 nrd=0.3 nrs=0.343056 sa=1.80167e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=19200 $Y=41510 $D=28
M3907 4033 4027 4032 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.85767e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=19680 $Y=41510 $D=28
M3908 4031 4030 4033 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10571e-13 as=1.08e-13 pd=9.71429e-07 ps=9.6e-07 nrd=0.307143 nrs=0.3 sa=1.91367e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=20160 $Y=41510 $D=28
M3909 VSS 4032 4031 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.63084e-13 as=1.21629e-13 pd=1.15677e-06 ps=1.06857e-06 nrd=0.374389 nrs=0.279221 sa=1.81515e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=20640 $Y=41450 $D=28
M3910 4032 94 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.27329e-13 pd=2.48e-06 ps=1.61247e-06 nrd=0.347826 nrs=0.268583 sa=1.46022e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=21200 $Y=41190 $D=28
M3911 VSS 4029 944 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=22160 $Y=41190 $D=28
M3912 8 4033 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=22640 $Y=41190 $D=28
M3913 4035 92 VSS VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.062e-13 as=1.888e-13 pd=9.5e-07 ps=1.82e-06 nrd=0.305085 nrs=0.542373 sa=3.2e-07 sb=1.14305e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=22010 $Y=48560 $D=28
M3914 VSS 92 4035 VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22021e-13 as=1.062e-13 pd=1.28489e-06 ps=9.5e-07 nrd=0.350534 nrs=0.305085 sa=8e-07 sb=6.63051e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=22490 $Y=48560 $D=28
M3915 4034 92 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=9.92711e-14 pd=1.6e-06 ps=1.04533e-06 nrd=0.666667 nrs=0.430864 sa=1.24e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=22930 $Y=48670 $D=28
M3916 VSS 4034 4036 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47609e-13 as=1.696e-13 pd=1.16284e-06 ps=1.7e-06 nrd=0.525486 nrs=0.603774 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=23970 $Y=48620 $D=28
M3917 4036 4034 VSS VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.54e-14 as=1.47609e-13 pd=8.9e-07 ps=1.16284e-06 nrd=0.339623 nrs=0.525486 sa=8.8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=24530 $Y=48620 $D=28
M3918 4037 120 4036 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.34138e-13 as=9.54e-14 pd=1.07927e-06 ps=8.9e-07 nrd=0.47753 nrs=0.339623 sa=1.36e-06 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=25010 $Y=48620 $D=28
M3919 4036 120 4037 VSS lpnfet w=5.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.824e-13 as=1.44262e-13 pd=1.78e-06 ps=1.16073e-06 nrd=0.561404 nrs=0.444019 sa=1.81053e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=25570 $Y=48620 $D=28
M3920 4037 4038 4035 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=26510 $Y=48710 $D=28
M3921 4035 4038 4037 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=26990 $Y=48710 $D=28
M3922 4040 120 4035 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=27470 $Y=48710 $D=28
M3923 4035 120 4040 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=27950 $Y=48710 $D=28
M3924 4036 4038 4040 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21e-13 as=3.016e-13 pd=9.9e-07 ps=2.56e-06 nrd=0.4 nrs=0.997025 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=28990 $Y=48760 $D=28
M3925 4040 4038 4036 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.016e-13 as=1.21e-13 pd=2.56e-06 ps=9.9e-07 nrd=0.997025 nrs=0.4 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=29550 $Y=48760 $D=28
M3926 VSS 120 4038 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.18002e-13 as=3.464e-13 pd=1.3493e-06 ps=2.52e-06 nrd=0.377428 nrs=0.599723 sa=4.3e-07 sb=1.71605e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=30740 $Y=48480 $D=28
M3927 4038 120 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45741e-13 as=2.18002e-13 pd=1.25176e-06 ps=1.3493e-06 nrd=0.252322 nrs=0.377428 sa=1.09e-06 sb=1.51632e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=31400 $Y=48480 $D=28
M3928 4039 4037 4038 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.235e-13 as=1.15059e-13 pd=1.07e-06 ps=9.88235e-07 nrd=0.343056 nrs=0.319608 sa=1.57e-06 sb=1.79e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=31880 $Y=48640 $D=28
M3929 4042 4040 4039 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.235e-13 pd=9.6e-07 ps=1.07e-06 nrd=0.3 nrs=0.343056 sa=1.80167e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=32400 $Y=48710 $D=28
M3930 4043 4037 4042 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.85767e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=32880 $Y=48710 $D=28
M3931 4041 4040 4043 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10571e-13 as=1.08e-13 pd=9.71429e-07 ps=9.6e-07 nrd=0.307143 nrs=0.3 sa=1.91367e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=33360 $Y=48710 $D=28
M3932 VSS 4042 4041 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.63084e-13 as=1.21629e-13 pd=1.15677e-06 ps=1.06857e-06 nrd=0.374389 nrs=0.279221 sa=1.81515e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=33840 $Y=48650 $D=28
M3933 4042 197 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.27329e-13 pd=2.48e-06 ps=1.61247e-06 nrd=0.347826 nrs=0.268583 sa=1.46022e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=34400 $Y=48390 $D=28
M3934 VSS 4039 121 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=35360 $Y=48390 $D=28
M3935 124 4043 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=35840 $Y=48390 $D=28
M3936 4045 77 VSS VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.062e-13 as=1.888e-13 pd=9.5e-07 ps=1.82e-06 nrd=0.305085 nrs=0.542373 sa=3.2e-07 sb=1.14305e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=23610 $Y=25250 $D=28
M3937 VSS 77 4045 VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22021e-13 as=1.062e-13 pd=1.28489e-06 ps=9.5e-07 nrd=0.350534 nrs=0.305085 sa=8e-07 sb=6.63051e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=24090 $Y=25250 $D=28
M3938 4044 77 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=9.92711e-14 pd=1.6e-06 ps=1.04533e-06 nrd=0.666667 nrs=0.430864 sa=1.24e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=24530 $Y=25250 $D=28
M3939 VSS 4044 4046 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47609e-13 as=1.696e-13 pd=1.16284e-06 ps=1.7e-06 nrd=0.525486 nrs=0.603774 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=25570 $Y=25250 $D=28
M3940 4046 4044 VSS VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.54e-14 as=1.47609e-13 pd=8.9e-07 ps=1.16284e-06 nrd=0.339623 nrs=0.525486 sa=8.8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=26130 $Y=25250 $D=28
M3941 4047 155 4046 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.34138e-13 as=9.54e-14 pd=1.07927e-06 ps=8.9e-07 nrd=0.47753 nrs=0.339623 sa=1.36e-06 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=26610 $Y=25250 $D=28
M3942 4046 155 4047 VSS lpnfet w=5.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.824e-13 as=1.44262e-13 pd=1.78e-06 ps=1.16073e-06 nrd=0.561404 nrs=0.444019 sa=1.81053e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=27170 $Y=25210 $D=28
M3943 4047 4048 4045 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=28110 $Y=25140 $D=28
M3944 4045 4048 4047 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=28590 $Y=25140 $D=28
M3945 4050 155 4045 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=29070 $Y=25140 $D=28
M3946 4045 155 4050 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=29550 $Y=25140 $D=28
M3947 4046 4048 4050 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21e-13 as=3.016e-13 pd=9.9e-07 ps=2.56e-06 nrd=0.4 nrs=0.997025 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=30590 $Y=25090 $D=28
M3948 4050 4048 4046 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.016e-13 as=1.21e-13 pd=2.56e-06 ps=9.9e-07 nrd=0.997025 nrs=0.4 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=31150 $Y=25090 $D=28
M3949 VSS 155 4048 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.18002e-13 as=3.464e-13 pd=1.3493e-06 ps=2.52e-06 nrd=0.377428 nrs=0.599723 sa=4.3e-07 sb=1.71605e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=32340 $Y=25160 $D=28
M3950 4048 155 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45741e-13 as=2.18002e-13 pd=1.25176e-06 ps=1.3493e-06 nrd=0.252322 nrs=0.377428 sa=1.09e-06 sb=1.51632e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=33000 $Y=25160 $D=28
M3951 4049 4047 4048 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.235e-13 as=1.15059e-13 pd=1.07e-06 ps=9.88235e-07 nrd=0.343056 nrs=0.319608 sa=1.57e-06 sb=1.79e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=33480 $Y=25160 $D=28
M3952 4052 4050 4049 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.235e-13 pd=9.6e-07 ps=1.07e-06 nrd=0.3 nrs=0.343056 sa=1.80167e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=34000 $Y=25090 $D=28
M3953 4053 4047 4052 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.85767e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=34480 $Y=25090 $D=28
M3954 4051 4050 4053 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10571e-13 as=1.08e-13 pd=9.71429e-07 ps=9.6e-07 nrd=0.307143 nrs=0.3 sa=1.91367e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=34960 $Y=25090 $D=28
M3955 VSS 4052 4051 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.63084e-13 as=1.21629e-13 pd=1.15677e-06 ps=1.06857e-06 nrd=0.374389 nrs=0.279221 sa=1.81515e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=35440 $Y=25090 $D=28
M3956 4052 126 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.27329e-13 pd=2.48e-06 ps=1.61247e-06 nrd=0.347826 nrs=0.268583 sa=1.46022e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=36000 $Y=25090 $D=28
M3957 VSS 4049 133 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=36960 $Y=25090 $D=28
M3958 130 4053 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=37440 $Y=25090 $D=28
M3959 4055 149 VSS VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.062e-13 as=1.888e-13 pd=9.5e-07 ps=1.82e-06 nrd=0.305085 nrs=0.542373 sa=3.2e-07 sb=1.14305e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=38810 $Y=70160 $D=28
M3960 VSS 149 4055 VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22021e-13 as=1.062e-13 pd=1.28489e-06 ps=9.5e-07 nrd=0.350534 nrs=0.305085 sa=8e-07 sb=6.63051e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=39290 $Y=70160 $D=28
M3961 4054 149 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=9.92711e-14 pd=1.6e-06 ps=1.04533e-06 nrd=0.666667 nrs=0.430864 sa=1.24e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=39730 $Y=70270 $D=28
M3962 VSS 4054 4056 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47609e-13 as=1.696e-13 pd=1.16284e-06 ps=1.7e-06 nrd=0.525486 nrs=0.603774 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=40770 $Y=70220 $D=28
M3963 4056 4054 VSS VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.54e-14 as=1.47609e-13 pd=8.9e-07 ps=1.16284e-06 nrd=0.339623 nrs=0.525486 sa=8.8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=41330 $Y=70220 $D=28
M3964 4057 225 4056 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.34138e-13 as=9.54e-14 pd=1.07927e-06 ps=8.9e-07 nrd=0.47753 nrs=0.339623 sa=1.36e-06 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=41810 $Y=70220 $D=28
M3965 4056 225 4057 VSS lpnfet w=5.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.824e-13 as=1.44262e-13 pd=1.78e-06 ps=1.16073e-06 nrd=0.561404 nrs=0.444019 sa=1.81053e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=42370 $Y=70220 $D=28
M3966 4057 4058 4055 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=43310 $Y=70310 $D=28
M3967 4055 4058 4057 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=43790 $Y=70310 $D=28
M3968 4060 225 4055 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=44270 $Y=70310 $D=28
M3969 4055 225 4060 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=44750 $Y=70310 $D=28
M3970 4056 4058 4060 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21e-13 as=3.016e-13 pd=9.9e-07 ps=2.56e-06 nrd=0.4 nrs=0.997025 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=45790 $Y=70360 $D=28
M3971 4060 4058 4056 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.016e-13 as=1.21e-13 pd=2.56e-06 ps=9.9e-07 nrd=0.997025 nrs=0.4 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=46350 $Y=70360 $D=28
M3972 VSS 225 4058 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.18002e-13 as=3.464e-13 pd=1.3493e-06 ps=2.52e-06 nrd=0.377428 nrs=0.599723 sa=4.3e-07 sb=1.71605e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=47540 $Y=70080 $D=28
M3973 4058 225 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45741e-13 as=2.18002e-13 pd=1.25176e-06 ps=1.3493e-06 nrd=0.252322 nrs=0.377428 sa=1.09e-06 sb=1.51632e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=48200 $Y=70080 $D=28
M3974 4059 4057 4058 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.235e-13 as=1.15059e-13 pd=1.07e-06 ps=9.88235e-07 nrd=0.343056 nrs=0.319608 sa=1.57e-06 sb=1.79e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=48680 $Y=70240 $D=28
M3975 4062 4060 4059 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.235e-13 pd=9.6e-07 ps=1.07e-06 nrd=0.3 nrs=0.343056 sa=1.80167e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=49200 $Y=70310 $D=28
M3976 4063 4057 4062 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.85767e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=49680 $Y=70310 $D=28
M3977 4061 4060 4063 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10571e-13 as=1.08e-13 pd=9.71429e-07 ps=9.6e-07 nrd=0.307143 nrs=0.3 sa=1.91367e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=50160 $Y=70310 $D=28
M3978 VSS 4062 4061 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.63084e-13 as=1.21629e-13 pd=1.15677e-06 ps=1.06857e-06 nrd=0.374389 nrs=0.279221 sa=1.81515e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=50640 $Y=70250 $D=28
M3979 4062 196 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.27329e-13 pd=2.48e-06 ps=1.61247e-06 nrd=0.347826 nrs=0.268583 sa=1.46022e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=51200 $Y=69990 $D=28
M3980 VSS 4059 191 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=52160 $Y=69990 $D=28
M3981 69 4063 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=52640 $Y=69990 $D=28
M3982 4065 152 VSS VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.062e-13 as=1.888e-13 pd=9.5e-07 ps=1.82e-06 nrd=0.305085 nrs=0.542373 sa=3.2e-07 sb=1.14305e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=39210 $Y=68450 $D=28
M3983 VSS 152 4065 VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22021e-13 as=1.062e-13 pd=1.28489e-06 ps=9.5e-07 nrd=0.350534 nrs=0.305085 sa=8e-07 sb=6.63051e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=39690 $Y=68450 $D=28
M3984 4064 152 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=9.92711e-14 pd=1.6e-06 ps=1.04533e-06 nrd=0.666667 nrs=0.430864 sa=1.24e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=40130 $Y=68450 $D=28
M3985 VSS 4064 4066 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47609e-13 as=1.696e-13 pd=1.16284e-06 ps=1.7e-06 nrd=0.525486 nrs=0.603774 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=41170 $Y=68450 $D=28
M3986 4066 4064 VSS VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.54e-14 as=1.47609e-13 pd=8.9e-07 ps=1.16284e-06 nrd=0.339623 nrs=0.525486 sa=8.8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=41730 $Y=68450 $D=28
M3987 4067 250 4066 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.34138e-13 as=9.54e-14 pd=1.07927e-06 ps=8.9e-07 nrd=0.47753 nrs=0.339623 sa=1.36e-06 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=42210 $Y=68450 $D=28
M3988 4066 250 4067 VSS lpnfet w=5.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.824e-13 as=1.44262e-13 pd=1.78e-06 ps=1.16073e-06 nrd=0.561404 nrs=0.444019 sa=1.81053e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=42770 $Y=68410 $D=28
M3989 4067 4068 4065 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=43710 $Y=68340 $D=28
M3990 4065 4068 4067 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=44190 $Y=68340 $D=28
M3991 4070 250 4065 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=44670 $Y=68340 $D=28
M3992 4065 250 4070 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=45150 $Y=68340 $D=28
M3993 4066 4068 4070 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21e-13 as=3.016e-13 pd=9.9e-07 ps=2.56e-06 nrd=0.4 nrs=0.997025 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=46190 $Y=68290 $D=28
M3994 4070 4068 4066 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.016e-13 as=1.21e-13 pd=2.56e-06 ps=9.9e-07 nrd=0.997025 nrs=0.4 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=46750 $Y=68290 $D=28
M3995 VSS 250 4068 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.18002e-13 as=3.464e-13 pd=1.3493e-06 ps=2.52e-06 nrd=0.377428 nrs=0.599723 sa=4.3e-07 sb=1.71605e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=47940 $Y=68360 $D=28
M3996 4068 250 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45741e-13 as=2.18002e-13 pd=1.25176e-06 ps=1.3493e-06 nrd=0.252322 nrs=0.377428 sa=1.09e-06 sb=1.51632e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=48600 $Y=68360 $D=28
M3997 4069 4067 4068 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.235e-13 as=1.15059e-13 pd=1.07e-06 ps=9.88235e-07 nrd=0.343056 nrs=0.319608 sa=1.57e-06 sb=1.79e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=49080 $Y=68360 $D=28
M3998 4072 4070 4069 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.235e-13 pd=9.6e-07 ps=1.07e-06 nrd=0.3 nrs=0.343056 sa=1.80167e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=49600 $Y=68290 $D=28
M3999 4073 4067 4072 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.85767e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=50080 $Y=68290 $D=28
M4000 4071 4070 4073 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10571e-13 as=1.08e-13 pd=9.71429e-07 ps=9.6e-07 nrd=0.307143 nrs=0.3 sa=1.91367e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=50560 $Y=68290 $D=28
M4001 VSS 4072 4071 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.63084e-13 as=1.21629e-13 pd=1.15677e-06 ps=1.06857e-06 nrd=0.374389 nrs=0.279221 sa=1.81515e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=51040 $Y=68290 $D=28
M4002 4072 190 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.27329e-13 pd=2.48e-06 ps=1.61247e-06 nrd=0.347826 nrs=0.268583 sa=1.46022e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=51600 $Y=68290 $D=28
M4003 VSS 4069 268 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=52560 $Y=68290 $D=28
M4004 196 4073 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=53040 $Y=68290 $D=28
M4005 4075 279 VSS VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.062e-13 as=1.888e-13 pd=9.5e-07 ps=1.82e-06 nrd=0.305085 nrs=0.542373 sa=3.2e-07 sb=1.14305e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=40810 $Y=46850 $D=28
M4006 VSS 279 4075 VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22021e-13 as=1.062e-13 pd=1.28489e-06 ps=9.5e-07 nrd=0.350534 nrs=0.305085 sa=8e-07 sb=6.63051e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=41290 $Y=46850 $D=28
M4007 4074 279 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=9.92711e-14 pd=1.6e-06 ps=1.04533e-06 nrd=0.666667 nrs=0.430864 sa=1.24e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=41730 $Y=46850 $D=28
M4008 VSS 4074 4076 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47609e-13 as=1.696e-13 pd=1.16284e-06 ps=1.7e-06 nrd=0.525486 nrs=0.603774 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=42770 $Y=46850 $D=28
M4009 4076 4074 VSS VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.54e-14 as=1.47609e-13 pd=8.9e-07 ps=1.16284e-06 nrd=0.339623 nrs=0.525486 sa=8.8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=43330 $Y=46850 $D=28
M4010 4077 812 4076 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.34138e-13 as=9.54e-14 pd=1.07927e-06 ps=8.9e-07 nrd=0.47753 nrs=0.339623 sa=1.36e-06 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=43810 $Y=46850 $D=28
M4011 4076 812 4077 VSS lpnfet w=5.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.824e-13 as=1.44262e-13 pd=1.78e-06 ps=1.16073e-06 nrd=0.561404 nrs=0.444019 sa=1.81053e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=44370 $Y=46810 $D=28
M4012 4077 4078 4075 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=45310 $Y=46740 $D=28
M4013 4075 4078 4077 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=45790 $Y=46740 $D=28
M4014 4080 812 4075 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=46270 $Y=46740 $D=28
M4015 4075 812 4080 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=46750 $Y=46740 $D=28
M4016 4076 4078 4080 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21e-13 as=3.016e-13 pd=9.9e-07 ps=2.56e-06 nrd=0.4 nrs=0.997025 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=47790 $Y=46690 $D=28
M4017 4080 4078 4076 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.016e-13 as=1.21e-13 pd=2.56e-06 ps=9.9e-07 nrd=0.997025 nrs=0.4 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=48350 $Y=46690 $D=28
M4018 VSS 812 4078 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.18002e-13 as=3.464e-13 pd=1.3493e-06 ps=2.52e-06 nrd=0.377428 nrs=0.599723 sa=4.3e-07 sb=1.71605e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=49540 $Y=46760 $D=28
M4019 4078 812 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45741e-13 as=2.18002e-13 pd=1.25176e-06 ps=1.3493e-06 nrd=0.252322 nrs=0.377428 sa=1.09e-06 sb=1.51632e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=50200 $Y=46760 $D=28
M4020 4079 4077 4078 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.235e-13 as=1.15059e-13 pd=1.07e-06 ps=9.88235e-07 nrd=0.343056 nrs=0.319608 sa=1.57e-06 sb=1.79e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=50680 $Y=46760 $D=28
M4021 4082 4080 4079 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.235e-13 pd=9.6e-07 ps=1.07e-06 nrd=0.3 nrs=0.343056 sa=1.80167e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=51200 $Y=46690 $D=28
M4022 4083 4077 4082 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.85767e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=51680 $Y=46690 $D=28
M4023 4081 4080 4083 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10571e-13 as=1.08e-13 pd=9.71429e-07 ps=9.6e-07 nrd=0.307143 nrs=0.3 sa=1.91367e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=52160 $Y=46690 $D=28
M4024 VSS 4082 4081 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.63084e-13 as=1.21629e-13 pd=1.15677e-06 ps=1.06857e-06 nrd=0.374389 nrs=0.279221 sa=1.81515e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=52640 $Y=46690 $D=28
M4025 4082 223 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.27329e-13 pd=2.48e-06 ps=1.61247e-06 nrd=0.347826 nrs=0.268583 sa=1.46022e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=53200 $Y=46690 $D=28
M4026 VSS 4079 149 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=54160 $Y=46690 $D=28
M4027 197 4083 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=54640 $Y=46690 $D=28
M4028 4085 331 VSS VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.062e-13 as=1.888e-13 pd=9.5e-07 ps=1.82e-06 nrd=0.305085 nrs=0.542373 sa=3.2e-07 sb=1.14305e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=84010 $Y=48560 $D=28
M4029 VSS 331 4085 VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22021e-13 as=1.062e-13 pd=1.28489e-06 ps=9.5e-07 nrd=0.350534 nrs=0.305085 sa=8e-07 sb=6.63051e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=84490 $Y=48560 $D=28
M4030 4084 331 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=9.92711e-14 pd=1.6e-06 ps=1.04533e-06 nrd=0.666667 nrs=0.430864 sa=1.24e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=84930 $Y=48670 $D=28
M4031 VSS 4084 4086 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47609e-13 as=1.696e-13 pd=1.16284e-06 ps=1.7e-06 nrd=0.525486 nrs=0.603774 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=85970 $Y=48620 $D=28
M4032 4086 4084 VSS VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.54e-14 as=1.47609e-13 pd=8.9e-07 ps=1.16284e-06 nrd=0.339623 nrs=0.525486 sa=8.8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=86530 $Y=48620 $D=28
M4033 4087 340 4086 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.34138e-13 as=9.54e-14 pd=1.07927e-06 ps=8.9e-07 nrd=0.47753 nrs=0.339623 sa=1.36e-06 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=87010 $Y=48620 $D=28
M4034 4086 340 4087 VSS lpnfet w=5.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.824e-13 as=1.44262e-13 pd=1.78e-06 ps=1.16073e-06 nrd=0.561404 nrs=0.444019 sa=1.81053e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=87570 $Y=48620 $D=28
M4035 4087 4088 4085 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=88510 $Y=48710 $D=28
M4036 4085 4088 4087 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=88990 $Y=48710 $D=28
M4037 4090 340 4085 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=89470 $Y=48710 $D=28
M4038 4085 340 4090 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=89950 $Y=48710 $D=28
M4039 4086 4088 4090 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21e-13 as=3.016e-13 pd=9.9e-07 ps=2.56e-06 nrd=0.4 nrs=0.997025 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=90990 $Y=48760 $D=28
M4040 4090 4088 4086 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.016e-13 as=1.21e-13 pd=2.56e-06 ps=9.9e-07 nrd=0.997025 nrs=0.4 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=91550 $Y=48760 $D=28
M4041 VSS 340 4088 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.18002e-13 as=3.464e-13 pd=1.3493e-06 ps=2.52e-06 nrd=0.377428 nrs=0.599723 sa=4.3e-07 sb=1.71605e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=92740 $Y=48480 $D=28
M4042 4088 340 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45741e-13 as=2.18002e-13 pd=1.25176e-06 ps=1.3493e-06 nrd=0.252322 nrs=0.377428 sa=1.09e-06 sb=1.51632e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=93400 $Y=48480 $D=28
M4043 4089 4087 4088 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.235e-13 as=1.15059e-13 pd=1.07e-06 ps=9.88235e-07 nrd=0.343056 nrs=0.319608 sa=1.57e-06 sb=1.79e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=93880 $Y=48640 $D=28
M4044 4092 4090 4089 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.235e-13 pd=9.6e-07 ps=1.07e-06 nrd=0.3 nrs=0.343056 sa=1.80167e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=94400 $Y=48710 $D=28
M4045 4093 4087 4092 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.85767e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=94880 $Y=48710 $D=28
M4046 4091 4090 4093 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10571e-13 as=1.08e-13 pd=9.71429e-07 ps=9.6e-07 nrd=0.307143 nrs=0.3 sa=1.91367e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=95360 $Y=48710 $D=28
M4047 VSS 4092 4091 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.63084e-13 as=1.21629e-13 pd=1.15677e-06 ps=1.06857e-06 nrd=0.374389 nrs=0.279221 sa=1.81515e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=95840 $Y=48650 $D=28
M4048 4092 355 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.27329e-13 pd=2.48e-06 ps=1.61247e-06 nrd=0.347826 nrs=0.268583 sa=1.46022e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=96400 $Y=48390 $D=28
M4049 VSS 4089 381 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=97360 $Y=48390 $D=28
M4050 831 4093 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=97840 $Y=48390 $D=28
M4051 4095 452 VSS VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.062e-13 as=1.888e-13 pd=9.5e-07 ps=1.82e-06 nrd=0.305085 nrs=0.542373 sa=3.2e-07 sb=1.14305e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=106810 $Y=34160 $D=28
M4052 VSS 452 4095 VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22021e-13 as=1.062e-13 pd=1.28489e-06 ps=9.5e-07 nrd=0.350534 nrs=0.305085 sa=8e-07 sb=6.63051e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=107290 $Y=34160 $D=28
M4053 4094 452 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=9.92711e-14 pd=1.6e-06 ps=1.04533e-06 nrd=0.666667 nrs=0.430864 sa=1.24e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=107730 $Y=34270 $D=28
M4054 VSS 4094 4096 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47609e-13 as=1.696e-13 pd=1.16284e-06 ps=1.7e-06 nrd=0.525486 nrs=0.603774 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=108770 $Y=34220 $D=28
M4055 4096 4094 VSS VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.54e-14 as=1.47609e-13 pd=8.9e-07 ps=1.16284e-06 nrd=0.339623 nrs=0.525486 sa=8.8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=109330 $Y=34220 $D=28
M4056 4097 418 4096 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.34138e-13 as=9.54e-14 pd=1.07927e-06 ps=8.9e-07 nrd=0.47753 nrs=0.339623 sa=1.36e-06 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=109810 $Y=34220 $D=28
M4057 4096 418 4097 VSS lpnfet w=5.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.824e-13 as=1.44262e-13 pd=1.78e-06 ps=1.16073e-06 nrd=0.561404 nrs=0.444019 sa=1.81053e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=110370 $Y=34220 $D=28
M4058 4097 4098 4095 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=111310 $Y=34310 $D=28
M4059 4095 4098 4097 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=111790 $Y=34310 $D=28
M4060 4100 418 4095 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=112270 $Y=34310 $D=28
M4061 4095 418 4100 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=112750 $Y=34310 $D=28
M4062 4096 4098 4100 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21e-13 as=3.016e-13 pd=9.9e-07 ps=2.56e-06 nrd=0.4 nrs=0.997025 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=113790 $Y=34360 $D=28
M4063 4100 4098 4096 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.016e-13 as=1.21e-13 pd=2.56e-06 ps=9.9e-07 nrd=0.997025 nrs=0.4 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=114350 $Y=34360 $D=28
M4064 VSS 418 4098 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.18002e-13 as=3.464e-13 pd=1.3493e-06 ps=2.52e-06 nrd=0.377428 nrs=0.599723 sa=4.3e-07 sb=1.71605e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=115540 $Y=34080 $D=28
M4065 4098 418 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45741e-13 as=2.18002e-13 pd=1.25176e-06 ps=1.3493e-06 nrd=0.252322 nrs=0.377428 sa=1.09e-06 sb=1.51632e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=116200 $Y=34080 $D=28
M4066 4099 4097 4098 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.235e-13 as=1.15059e-13 pd=1.07e-06 ps=9.88235e-07 nrd=0.343056 nrs=0.319608 sa=1.57e-06 sb=1.79e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=116680 $Y=34240 $D=28
M4067 4102 4100 4099 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.235e-13 pd=9.6e-07 ps=1.07e-06 nrd=0.3 nrs=0.343056 sa=1.80167e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=117200 $Y=34310 $D=28
M4068 4103 4097 4102 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.85767e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=117680 $Y=34310 $D=28
M4069 4101 4100 4103 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10571e-13 as=1.08e-13 pd=9.71429e-07 ps=9.6e-07 nrd=0.307143 nrs=0.3 sa=1.91367e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=118160 $Y=34310 $D=28
M4070 VSS 4102 4101 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.63084e-13 as=1.21629e-13 pd=1.15677e-06 ps=1.06857e-06 nrd=0.374389 nrs=0.279221 sa=1.81515e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=118640 $Y=34250 $D=28
M4071 4102 446 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.27329e-13 pd=2.48e-06 ps=1.61247e-06 nrd=0.347826 nrs=0.268583 sa=1.46022e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=119200 $Y=33990 $D=28
M4072 VSS 4099 451 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=120160 $Y=33990 $D=28
M4073 455 4103 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=120640 $Y=33990 $D=28
M4074 4105 413 VSS VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.062e-13 as=1.888e-13 pd=9.5e-07 ps=1.82e-06 nrd=0.305085 nrs=0.542373 sa=3.2e-07 sb=1.14305e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=110810 $Y=26960 $D=28
M4075 VSS 413 4105 VSS lpnfet w=5.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22021e-13 as=1.062e-13 pd=1.28489e-06 ps=9.5e-07 nrd=0.350534 nrs=0.305085 sa=8e-07 sb=6.63051e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=111290 $Y=26960 $D=28
M4076 4104 413 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.536e-13 as=9.92711e-14 pd=1.6e-06 ps=1.04533e-06 nrd=0.666667 nrs=0.430864 sa=1.24e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=111730 $Y=27070 $D=28
M4077 VSS 4104 4106 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.47609e-13 as=1.696e-13 pd=1.16284e-06 ps=1.7e-06 nrd=0.525486 nrs=0.603774 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=112770 $Y=27020 $D=28
M4078 4106 4104 VSS VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.54e-14 as=1.47609e-13 pd=8.9e-07 ps=1.16284e-06 nrd=0.339623 nrs=0.525486 sa=8.8e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=113330 $Y=27020 $D=28
M4079 4107 455 4106 VSS lpnfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.34138e-13 as=9.54e-14 pd=1.07927e-06 ps=8.9e-07 nrd=0.47753 nrs=0.339623 sa=1.36e-06 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=113810 $Y=27020 $D=28
M4080 4106 455 4107 VSS lpnfet w=5.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.824e-13 as=1.44262e-13 pd=1.78e-06 ps=1.16073e-06 nrd=0.561404 nrs=0.444019 sa=1.81053e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.28e-14 panw9=0 panw10=0 $X=114370 $Y=27020 $D=28
M4081 4107 4108 4105 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=115310 $Y=27110 $D=28
M4082 4105 4108 4107 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=115790 $Y=27110 $D=28
M4083 4110 455 4105 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=9.9e-14 pd=9.1e-07 ps=9.1e-07 nrd=0.327273 nrs=0.327273 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=116270 $Y=27110 $D=28
M4084 4105 455 4110 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76e-13 as=9.9e-14 pd=1.74e-06 ps=9.1e-07 nrd=0.581818 nrs=0.327273 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=116750 $Y=27110 $D=28
M4085 4106 4108 4110 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21e-13 as=3.016e-13 pd=9.9e-07 ps=2.56e-06 nrd=0.4 nrs=0.997025 sa=3.6e-07 sb=9.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=117790 $Y=27160 $D=28
M4086 4110 4108 4106 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.016e-13 as=1.21e-13 pd=2.56e-06 ps=9.9e-07 nrd=0.997025 nrs=0.4 sa=9.2e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=118350 $Y=27160 $D=28
M4087 VSS 455 4108 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.18002e-13 as=3.464e-13 pd=1.3493e-06 ps=2.52e-06 nrd=0.377428 nrs=0.599723 sa=4.3e-07 sb=1.71605e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=119540 $Y=26880 $D=28
M4088 4108 455 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45741e-13 as=2.18002e-13 pd=1.25176e-06 ps=1.3493e-06 nrd=0.252322 nrs=0.377428 sa=1.09e-06 sb=1.51632e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=120200 $Y=26880 $D=28
M4089 4109 4107 4108 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.235e-13 as=1.15059e-13 pd=1.07e-06 ps=9.88235e-07 nrd=0.343056 nrs=0.319608 sa=1.57e-06 sb=1.79e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=120680 $Y=27040 $D=28
M4090 4112 4110 4109 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.235e-13 pd=9.6e-07 ps=1.07e-06 nrd=0.3 nrs=0.343056 sa=1.80167e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=121200 $Y=27110 $D=28
M4091 4113 4107 4112 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.85767e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=121680 $Y=27110 $D=28
M4092 4111 4110 4113 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10571e-13 as=1.08e-13 pd=9.71429e-07 ps=9.6e-07 nrd=0.307143 nrs=0.3 sa=1.91367e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=122160 $Y=27110 $D=28
M4093 VSS 4112 4111 VSS lpnfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.63084e-13 as=1.21629e-13 pd=1.15677e-06 ps=1.06857e-06 nrd=0.374389 nrs=0.279221 sa=1.81515e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=122640 $Y=27050 $D=28
M4094 4112 461 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.27329e-13 pd=2.48e-06 ps=1.61247e-06 nrd=0.347826 nrs=0.268583 sa=1.46022e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=123200 $Y=26790 $D=28
M4095 VSS 4109 463 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=124160 $Y=26790 $D=28
M4096 448 4113 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.128e-13 as=1.656e-13 pd=2.52e-06 ps=1.28e-06 nrd=0.369565 nrs=0.195652 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=124640 $Y=26790 $D=28
M4097 VSS 30 4114 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.26304e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=16860 $Y=48390 $D=28
M4098 4114 43 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=8e-07 sb=7.83043e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=17340 $Y=48390 $D=28
M4099 4115 61 4114 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.788e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.329395 nrs=0.195652 sa=1.28e-06 sb=3.03043e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=17820 $Y=48390 $D=28
M4100 75 4115 VSS VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46824e-13 as=2.496e-13 pd=1.17459e-06 ps=2.2e-06 nrd=0.241327 nrs=0.410256 sa=3.2e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=18780 $Y=48530 $D=28
M4101 VSS 4115 75 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.73176e-13 pd=2.37667e-06 ps=1.38541e-06 nrd=0.368478 nrs=0.204604 sa=7.2087e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=19260 $Y=48390 $D=28
M4102 VSS 431 4117 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=1.26304e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=109660 $Y=75490 $D=28
M4103 4117 402 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=8e-07 sb=7.83043e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=110140 $Y=75490 $D=28
M4104 4118 435 4117 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.788e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.329395 nrs=0.195652 sa=1.28e-06 sb=3.03043e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=110620 $Y=75490 $D=28
M4105 415 4118 VSS VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46824e-13 as=2.496e-13 pd=1.17459e-06 ps=2.2e-06 nrd=0.241327 nrs=0.410256 sa=3.2e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=111580 $Y=75490 $D=28
M4106 VSS 4118 415 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.1188e-13 as=1.73176e-13 pd=2.37667e-06 ps=1.38541e-06 nrd=0.368478 nrs=0.204604 sa=7.2087e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=112060 $Y=75490 $D=28
M4107 VSS 74 4120 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.2973e-13 as=1.92e-13 pd=1.32162e-06 ps=1.84e-06 nrd=0.36036 nrs=0.533333 sa=3.2e-07 sb=1.72e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=23670 $Y=27110 $D=28
M4108 4120 57 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.2973e-13 pd=9.6e-07 ps=1.32162e-06 nrd=0.3 nrs=0.36036 sa=7.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=24110 $Y=27110 $D=28
M4109 77 84 4120 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.24e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=24590 $Y=27110 $D=28
M4110 4120 83 77 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.72e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=25070 $Y=27110 $D=28
M4111 VSS 102 4123 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.2973e-13 as=1.92e-13 pd=1.32162e-06 ps=1.84e-06 nrd=0.36036 nrs=0.533333 sa=3.2e-07 sb=1.72e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=29670 $Y=32290 $D=28
M4112 4123 74 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.2973e-13 pd=9.6e-07 ps=1.32162e-06 nrd=0.3 nrs=0.36036 sa=7.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=30110 $Y=32290 $D=28
M4113 106 84 4123 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.24e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=30590 $Y=32290 $D=28
M4114 4123 112 106 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.72e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=31070 $Y=32290 $D=28
M4115 VSS 148 4126 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.2973e-13 as=1.92e-13 pd=1.32162e-06 ps=1.84e-06 nrd=0.36036 nrs=0.533333 sa=3.2e-07 sb=1.72e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=38470 $Y=25090 $D=28
M4116 4126 144 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.2973e-13 pd=9.6e-07 ps=1.32162e-06 nrd=0.3 nrs=0.36036 sa=7.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=38910 $Y=25090 $D=28
M4117 155 182 4126 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.24e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=39390 $Y=25090 $D=28
M4118 4126 165 155 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.72e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=39870 $Y=25090 $D=28
M4119 VSS 148 4129 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.2973e-13 as=1.92e-13 pd=1.32162e-06 ps=1.84e-06 nrd=0.36036 nrs=0.533333 sa=3.2e-07 sb=1.72e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=40070 $Y=48710 $D=28
M4120 4129 166 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.2973e-13 pd=9.6e-07 ps=1.32162e-06 nrd=0.3 nrs=0.36036 sa=7.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=40510 $Y=48710 $D=28
M4121 178 164 4129 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.24e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=40990 $Y=48710 $D=28
M4122 4129 198 178 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.72e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=41470 $Y=48710 $D=28
M4123 VSS 148 4132 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.2973e-13 as=1.92e-13 pd=1.32162e-06 ps=1.84e-06 nrd=0.36036 nrs=0.533333 sa=3.2e-07 sb=1.72e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=42470 $Y=34310 $D=28
M4124 4132 164 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.2973e-13 pd=9.6e-07 ps=1.32162e-06 nrd=0.3 nrs=0.36036 sa=7.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=42910 $Y=34310 $D=28
M4125 93 198 4132 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.24e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=43390 $Y=34310 $D=28
M4126 4132 144 93 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.72e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=43870 $Y=34310 $D=28
M4127 VSS 293 4135 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.2973e-13 as=1.92e-13 pd=1.32162e-06 ps=1.84e-06 nrd=0.36036 nrs=0.533333 sa=3.2e-07 sb=1.72e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=73270 $Y=55910 $D=28
M4128 4135 325 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.2973e-13 pd=9.6e-07 ps=1.32162e-06 nrd=0.3 nrs=0.36036 sa=7.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=73710 $Y=55910 $D=28
M4129 288 295 4135 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.24e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=74190 $Y=55910 $D=28
M4130 4135 280 288 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.72e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=74670 $Y=55910 $D=28
M4131 VSS 343 4138 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.2973e-13 as=1.92e-13 pd=1.32162e-06 ps=1.84e-06 nrd=0.36036 nrs=0.533333 sa=3.2e-07 sb=1.72e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=88470 $Y=53890 $D=28
M4132 4138 325 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.2973e-13 pd=9.6e-07 ps=1.32162e-06 nrd=0.3 nrs=0.36036 sa=7.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=88910 $Y=53890 $D=28
M4133 331 295 4138 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.24e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=89390 $Y=53890 $D=28
M4134 4138 328 331 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.72e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=89870 $Y=53890 $D=28
M4135 VSS 400 4141 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.2973e-13 as=1.92e-13 pd=1.32162e-06 ps=1.84e-06 nrd=0.36036 nrs=0.533333 sa=3.2e-07 sb=1.72e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=108070 $Y=46690 $D=28
M4136 4141 406 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.2973e-13 pd=9.6e-07 ps=1.32162e-06 nrd=0.3 nrs=0.36036 sa=7.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=108510 $Y=46690 $D=28
M4137 910 416 4141 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.08e-13 as=1.08e-13 pd=9.6e-07 ps=9.6e-07 nrd=0.3 nrs=0.3 sa=1.24e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=108990 $Y=46690 $D=28
M4138 4141 410 910 VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92e-13 as=1.08e-13 pd=1.84e-06 ps=9.6e-07 nrd=0.533333 nrs=0.3 sa=1.72e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=109470 $Y=46690 $D=28
M4139 VSS 84 4144 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21101e-13 as=2.048e-13 pd=1.02582e-06 ps=1.92e-06 nrd=0.295656 nrs=0.5 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=17320 $Y=34270 $D=28
M4140 4144 57 VSS VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.45699e-13 pd=1.13e-06 ps=1.23418e-06 nrd=0.233766 nrs=0.24574 sa=7.12208e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=17800 $Y=34140 $D=28
M4141 VSS 57 4144 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44594e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.243876 nrs=0.233766 sa=1.19221e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=18280 $Y=34140 $D=28
M4142 4144 84 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.69006e-13 pd=1.26e-06 ps=1.35808e-06 nrd=0.2 nrs=0.208649 sa=1.47111e-06 sb=1.95956e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=18760 $Y=34010 $D=28
M4143 VSS 84 4144 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.78044e-06 sb=1.89022e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=19240 $Y=34010 $D=28
M4144 4144 57 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.89022e-06 sb=1.82089e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=19720 $Y=34010 $D=28
M4145 70 142 4144 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69006e-13 as=1.62e-13 pd=1.35808e-06 ps=1.26e-06 nrd=0.208649 nrs=0.2 sa=1.95956e-06 sb=1.75156e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=20200 $Y=34010 $D=28
M4146 4144 74 70 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.44594e-13 pd=1.13e-06 ps=1.16192e-06 nrd=0.233766 nrs=0.243876 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=20680 $Y=34140 $D=28
M4147 70 74 4144 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=21160 $Y=34140 $D=28
M4148 4144 142 70 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=21640 $Y=34140 $D=28
M4149 70 142 4144 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.40998e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.23781 nrs=0.233766 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=22120 $Y=34140 $D=28
M4150 4144 74 70 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.88e-13 as=1.64802e-13 pd=2.44e-06 ps=1.35808e-06 nrd=0.355556 nrs=0.20346 sa=1.74289e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=22600 $Y=34010 $D=28
M4151 VSS 181 4151 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21101e-13 as=2.048e-13 pd=1.02582e-06 ps=1.92e-06 nrd=0.295656 nrs=0.5 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=44520 $Y=61090 $D=28
M4152 4151 189 VSS VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.45699e-13 pd=1.13e-06 ps=1.23418e-06 nrd=0.233766 nrs=0.24574 sa=7.12208e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=45000 $Y=61090 $D=28
M4153 VSS 189 4151 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44594e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.243876 nrs=0.233766 sa=1.19221e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=45480 $Y=61090 $D=28
M4154 4151 181 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.69006e-13 pd=1.26e-06 ps=1.35808e-06 nrd=0.2 nrs=0.208649 sa=1.47111e-06 sb=1.95956e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=45960 $Y=61090 $D=28
M4155 VSS 181 4151 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.78044e-06 sb=1.89022e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=46440 $Y=61090 $D=28
M4156 4151 189 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.89022e-06 sb=1.82089e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=46920 $Y=61090 $D=28
M4157 273 179 4151 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69006e-13 as=1.62e-13 pd=1.35808e-06 ps=1.26e-06 nrd=0.208649 nrs=0.2 sa=1.95956e-06 sb=1.75156e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=47400 $Y=61090 $D=28
M4158 4151 151 273 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.44594e-13 pd=1.13e-06 ps=1.16192e-06 nrd=0.233766 nrs=0.243876 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=47880 $Y=61090 $D=28
M4159 273 151 4151 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=48360 $Y=61090 $D=28
M4160 4151 179 273 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=48840 $Y=61090 $D=28
M4161 273 179 4151 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.40998e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.23781 nrs=0.233766 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=49320 $Y=61090 $D=28
M4162 4151 151 273 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.88e-13 as=1.64802e-13 pd=2.44e-06 ps=1.35808e-06 nrd=0.355556 nrs=0.20346 sa=1.74289e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=49800 $Y=61090 $D=28
M4163 VSS 212 4158 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21101e-13 as=2.048e-13 pd=1.02582e-06 ps=1.92e-06 nrd=0.295656 nrs=0.5 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=52520 $Y=39490 $D=28
M4164 4158 199 VSS VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.45699e-13 pd=1.13e-06 ps=1.23418e-06 nrd=0.233766 nrs=0.24574 sa=7.12208e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=53000 $Y=39490 $D=28
M4165 VSS 199 4158 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44594e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.243876 nrs=0.233766 sa=1.19221e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=53480 $Y=39490 $D=28
M4166 4158 212 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.69006e-13 pd=1.26e-06 ps=1.35808e-06 nrd=0.2 nrs=0.208649 sa=1.47111e-06 sb=1.95956e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=53960 $Y=39490 $D=28
M4167 VSS 212 4158 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.78044e-06 sb=1.89022e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=54440 $Y=39490 $D=28
M4168 4158 199 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.89022e-06 sb=1.82089e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=54920 $Y=39490 $D=28
M4169 194 219 4158 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69006e-13 as=1.62e-13 pd=1.35808e-06 ps=1.26e-06 nrd=0.208649 nrs=0.2 sa=1.95956e-06 sb=1.75156e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=55400 $Y=39490 $D=28
M4170 4158 232 194 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.44594e-13 pd=1.13e-06 ps=1.16192e-06 nrd=0.233766 nrs=0.243876 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=55880 $Y=39490 $D=28
M4171 194 232 4158 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=56360 $Y=39490 $D=28
M4172 4158 219 194 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=56840 $Y=39490 $D=28
M4173 194 219 4158 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.40998e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.23781 nrs=0.233766 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=57320 $Y=39490 $D=28
M4174 4158 232 194 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.88e-13 as=1.64802e-13 pd=2.44e-06 ps=1.35808e-06 nrd=0.355556 nrs=0.20346 sa=1.74289e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=57800 $Y=39490 $D=28
M4175 VSS 199 4165 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21101e-13 as=2.048e-13 pd=1.02582e-06 ps=1.92e-06 nrd=0.295656 nrs=0.5 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=60920 $Y=34270 $D=28
M4176 4165 209 VSS VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.45699e-13 pd=1.13e-06 ps=1.23418e-06 nrd=0.233766 nrs=0.24574 sa=7.12208e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=61400 $Y=34140 $D=28
M4177 VSS 209 4165 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44594e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.243876 nrs=0.233766 sa=1.19221e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=61880 $Y=34140 $D=28
M4178 4165 199 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.69006e-13 pd=1.26e-06 ps=1.35808e-06 nrd=0.2 nrs=0.208649 sa=1.47111e-06 sb=1.95956e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=62360 $Y=34010 $D=28
M4179 VSS 199 4165 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.78044e-06 sb=1.89022e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=62840 $Y=34010 $D=28
M4180 4165 209 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.89022e-06 sb=1.82089e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=63320 $Y=34010 $D=28
M4181 224 231 4165 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69006e-13 as=1.62e-13 pd=1.35808e-06 ps=1.26e-06 nrd=0.208649 nrs=0.2 sa=1.95956e-06 sb=1.75156e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=63800 $Y=34010 $D=28
M4182 4165 242 224 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.44594e-13 pd=1.13e-06 ps=1.16192e-06 nrd=0.233766 nrs=0.243876 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=64280 $Y=34140 $D=28
M4183 224 242 4165 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=64760 $Y=34140 $D=28
M4184 4165 231 224 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=65240 $Y=34140 $D=28
M4185 224 231 4165 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.40998e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.23781 nrs=0.233766 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=65720 $Y=34140 $D=28
M4186 4165 242 224 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.88e-13 as=1.64802e-13 pd=2.44e-06 ps=1.35808e-06 nrd=0.355556 nrs=0.20346 sa=1.74289e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=66200 $Y=34010 $D=28
M4187 VSS 301 4172 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21101e-13 as=2.048e-13 pd=1.02582e-06 ps=1.92e-06 nrd=0.295656 nrs=0.5 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=69320 $Y=39490 $D=28
M4188 4172 267 VSS VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.45699e-13 pd=1.13e-06 ps=1.23418e-06 nrd=0.233766 nrs=0.24574 sa=7.12208e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=69800 $Y=39490 $D=28
M4189 VSS 267 4172 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44594e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.243876 nrs=0.233766 sa=1.19221e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=70280 $Y=39490 $D=28
M4190 4172 301 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.69006e-13 pd=1.26e-06 ps=1.35808e-06 nrd=0.2 nrs=0.208649 sa=1.47111e-06 sb=1.95956e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=70760 $Y=39490 $D=28
M4191 VSS 301 4172 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.78044e-06 sb=1.89022e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=71240 $Y=39490 $D=28
M4192 4172 267 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.89022e-06 sb=1.82089e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=71720 $Y=39490 $D=28
M4193 279 212 4172 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69006e-13 as=1.62e-13 pd=1.35808e-06 ps=1.26e-06 nrd=0.208649 nrs=0.2 sa=1.95956e-06 sb=1.75156e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=72200 $Y=39490 $D=28
M4194 4172 282 279 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.44594e-13 pd=1.13e-06 ps=1.16192e-06 nrd=0.233766 nrs=0.243876 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=72680 $Y=39490 $D=28
M4195 279 282 4172 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=73160 $Y=39490 $D=28
M4196 4172 212 279 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=73640 $Y=39490 $D=28
M4197 279 212 4172 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.40998e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.23781 nrs=0.233766 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=74120 $Y=39490 $D=28
M4198 4172 282 279 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.88e-13 as=1.64802e-13 pd=2.44e-06 ps=1.35808e-06 nrd=0.355556 nrs=0.20346 sa=1.74289e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=74600 $Y=39490 $D=28
M4199 VSS 328 4179 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21101e-13 as=2.048e-13 pd=1.02582e-06 ps=1.92e-06 nrd=0.295656 nrs=0.5 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=74520 $Y=48670 $D=28
M4200 4179 325 VSS VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.45699e-13 pd=1.13e-06 ps=1.23418e-06 nrd=0.233766 nrs=0.24574 sa=7.12208e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=75000 $Y=48540 $D=28
M4201 VSS 325 4179 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44594e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.243876 nrs=0.233766 sa=1.19221e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=75480 $Y=48540 $D=28
M4202 4179 328 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.69006e-13 pd=1.26e-06 ps=1.35808e-06 nrd=0.2 nrs=0.208649 sa=1.47111e-06 sb=1.95956e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=75960 $Y=48410 $D=28
M4203 VSS 328 4179 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.78044e-06 sb=1.89022e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=76440 $Y=48410 $D=28
M4204 4179 325 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.89022e-06 sb=1.82089e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=76920 $Y=48410 $D=28
M4205 341 293 4179 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69006e-13 as=1.62e-13 pd=1.35808e-06 ps=1.26e-06 nrd=0.208649 nrs=0.2 sa=1.95956e-06 sb=1.75156e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=77400 $Y=48410 $D=28
M4206 4179 295 341 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.44594e-13 pd=1.13e-06 ps=1.16192e-06 nrd=0.233766 nrs=0.243876 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=77880 $Y=48540 $D=28
M4207 341 295 4179 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=78360 $Y=48540 $D=28
M4208 4179 293 341 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=78840 $Y=48540 $D=28
M4209 341 293 4179 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.40998e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.23781 nrs=0.233766 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=79320 $Y=48540 $D=28
M4210 4179 295 341 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.88e-13 as=1.64802e-13 pd=2.44e-06 ps=1.35808e-06 nrd=0.355556 nrs=0.20346 sa=1.74289e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=79800 $Y=48410 $D=28
M4211 VSS 314 4186 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21101e-13 as=2.048e-13 pd=1.02582e-06 ps=1.92e-06 nrd=0.295656 nrs=0.5 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=89320 $Y=34270 $D=28
M4212 4186 336 VSS VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.45699e-13 pd=1.13e-06 ps=1.23418e-06 nrd=0.233766 nrs=0.24574 sa=7.12208e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=89800 $Y=34140 $D=28
M4213 VSS 336 4186 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44594e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.243876 nrs=0.233766 sa=1.19221e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=90280 $Y=34140 $D=28
M4214 4186 314 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.69006e-13 pd=1.26e-06 ps=1.35808e-06 nrd=0.2 nrs=0.208649 sa=1.47111e-06 sb=1.95956e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=90760 $Y=34010 $D=28
M4215 VSS 314 4186 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.78044e-06 sb=1.89022e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=91240 $Y=34010 $D=28
M4216 4186 336 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.89022e-06 sb=1.82089e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=91720 $Y=34010 $D=28
M4217 346 327 4186 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69006e-13 as=1.62e-13 pd=1.35808e-06 ps=1.26e-06 nrd=0.208649 nrs=0.2 sa=1.95956e-06 sb=1.75156e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=92200 $Y=34010 $D=28
M4218 4186 330 346 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.44594e-13 pd=1.13e-06 ps=1.16192e-06 nrd=0.233766 nrs=0.243876 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=92680 $Y=34140 $D=28
M4219 346 330 4186 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=93160 $Y=34140 $D=28
M4220 4186 327 346 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=93640 $Y=34140 $D=28
M4221 346 327 4186 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.40998e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.23781 nrs=0.233766 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=94120 $Y=34140 $D=28
M4222 4186 330 346 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.88e-13 as=1.64802e-13 pd=2.44e-06 ps=1.35808e-06 nrd=0.355556 nrs=0.20346 sa=1.74289e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=94600 $Y=34010 $D=28
M4223 VSS 336 4193 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21101e-13 as=2.048e-13 pd=1.02582e-06 ps=1.92e-06 nrd=0.295656 nrs=0.5 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=91720 $Y=41470 $D=28
M4224 4193 327 VSS VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.45699e-13 pd=1.13e-06 ps=1.23418e-06 nrd=0.233766 nrs=0.24574 sa=7.12208e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=92200 $Y=41340 $D=28
M4225 VSS 327 4193 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44594e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.243876 nrs=0.233766 sa=1.19221e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=92680 $Y=41340 $D=28
M4226 4193 336 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.69006e-13 pd=1.26e-06 ps=1.35808e-06 nrd=0.2 nrs=0.208649 sa=1.47111e-06 sb=1.95956e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=93160 $Y=41210 $D=28
M4227 VSS 336 4193 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.78044e-06 sb=1.89022e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=93640 $Y=41210 $D=28
M4228 4193 327 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.89022e-06 sb=1.82089e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=94120 $Y=41210 $D=28
M4229 348 319 4193 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69006e-13 as=1.62e-13 pd=1.35808e-06 ps=1.26e-06 nrd=0.208649 nrs=0.2 sa=1.95956e-06 sb=1.75156e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=94600 $Y=41210 $D=28
M4230 4193 330 348 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.44594e-13 pd=1.13e-06 ps=1.16192e-06 nrd=0.233766 nrs=0.243876 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=95080 $Y=41340 $D=28
M4231 348 330 4193 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=95560 $Y=41340 $D=28
M4232 4193 319 348 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=96040 $Y=41340 $D=28
M4233 348 319 4193 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.40998e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.23781 nrs=0.233766 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=96520 $Y=41340 $D=28
M4234 4193 330 348 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.88e-13 as=1.64802e-13 pd=2.44e-06 ps=1.35808e-06 nrd=0.355556 nrs=0.20346 sa=1.74289e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=97000 $Y=41210 $D=28
M4235 VSS 419 4200 VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.21101e-13 as=2.048e-13 pd=1.02582e-06 ps=1.92e-06 nrd=0.295656 nrs=0.5 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=107720 $Y=41470 $D=28
M4236 4200 400 VSS VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.45699e-13 pd=1.13e-06 ps=1.23418e-06 nrd=0.233766 nrs=0.24574 sa=7.12208e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=108200 $Y=41340 $D=28
M4237 VSS 400 4200 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44594e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.243876 nrs=0.233766 sa=1.19221e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=108680 $Y=41340 $D=28
M4238 4200 419 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.69006e-13 pd=1.26e-06 ps=1.35808e-06 nrd=0.2 nrs=0.208649 sa=1.47111e-06 sb=1.95956e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=109160 $Y=41210 $D=28
M4239 VSS 419 4200 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.78044e-06 sb=1.89022e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=109640 $Y=41210 $D=28
M4240 4200 400 VSS VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62e-13 as=1.62e-13 pd=1.26e-06 ps=1.26e-06 nrd=0.2 nrs=0.2 sa=1.89022e-06 sb=1.82089e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=110120 $Y=41210 $D=28
M4241 365 343 4200 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.69006e-13 as=1.62e-13 pd=1.35808e-06 ps=1.26e-06 nrd=0.208649 nrs=0.2 sa=1.95956e-06 sb=1.75156e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=110600 $Y=41210 $D=28
M4242 4200 410 365 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.44594e-13 pd=1.13e-06 ps=1.16192e-06 nrd=0.233766 nrs=0.243876 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=111080 $Y=41340 $D=28
M4243 365 410 4200 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=111560 $Y=41340 $D=28
M4244 4200 343 365 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=1.386e-13 pd=1.13e-06 ps=1.13e-06 nrd=0.233766 nrs=0.233766 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=112040 $Y=41340 $D=28
M4245 365 343 4200 VSS lpnfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.40998e-13 as=1.386e-13 pd=1.16192e-06 ps=1.13e-06 nrd=0.23781 nrs=0.233766 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=112520 $Y=41340 $D=28
M4246 4200 410 365 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.88e-13 as=1.64802e-13 pd=2.44e-06 ps=1.35808e-06 nrd=0.355556 nrs=0.20346 sa=1.74289e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=113000 $Y=41210 $D=28
M4247 4209 148 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.8e-14 as=2.25853e-13 pd=6.8e-07 ps=1.89474e-06 nrd=0.208333 nrs=0.980263 sa=3.6e-07 sb=1.5e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=53560 $Y=55980 $D=28
M4248 4208 168 4209 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.32571e-14 as=4.8e-14 pd=9.6e-07 ps=6.8e-07 nrd=0.404762 nrs=0.208333 sa=6.8e-07 sb=1.18e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=53880 $Y=55980 $D=28
M4249 VSS 200 4208 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30308e-13 as=6.99429e-14 pd=8.38033e-07 ps=7.2e-07 nrd=1.00546 nrs=0.539683 sa=1.16e-06 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=54360 $Y=56100 $D=28
M4250 234 4208 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.752e-13 as=3.11292e-13 pd=2.36e-06 ps=2.00197e-06 nrd=0.372093 nrs=0.420892 sa=1.0493e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=55040 $Y=55600 $D=28
M4251 4212 400 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.8e-14 as=2.25853e-13 pd=6.8e-07 ps=1.89474e-06 nrd=0.208333 nrs=0.980263 sa=3.6e-07 sb=1.5e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=105560 $Y=46740 $D=28
M4252 4211 410 4212 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.32571e-14 as=4.8e-14 pd=9.6e-07 ps=6.8e-07 nrd=0.404762 nrs=0.208333 sa=6.8e-07 sb=1.18e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=105880 $Y=46740 $D=28
M4253 VSS 406 4211 VSS lpnfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30308e-13 as=6.99429e-14 pd=8.38033e-07 ps=7.2e-07 nrd=1.00546 nrs=0.539683 sa=1.16e-06 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=106360 $Y=46740 $D=28
M4254 403 4211 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.752e-13 as=3.11292e-13 pd=2.36e-06 ps=2.00197e-06 nrd=0.372093 nrs=0.420892 sa=1.0493e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=107040 $Y=46740 $D=28
M4255 110 89 VSS VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.46e-14 as=1.99029e-13 pd=8.3e-07 ps=1.70453e-06 nrd=0.382979 nrs=0.900993 sa=3.6e-07 sb=8.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=32900 $Y=63050 $D=28
M4256 VSS 89 110 VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.927e-13 as=8.46e-14 pd=1.76e-06 ps=8.3e-07 nrd=0.87234 nrs=0.382979 sa=8.4e-07 sb=4.1e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=33380 $Y=63050 $D=28
M4257 371 344 VSS VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.46e-14 as=1.99029e-13 pd=8.3e-07 ps=1.70453e-06 nrd=0.382979 nrs=0.900993 sa=3.6e-07 sb=8.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=100900 $Y=12650 $D=28
M4258 VSS 344 371 VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.927e-13 as=8.46e-14 pd=1.76e-06 ps=8.3e-07 nrd=0.87234 nrs=0.382979 sa=8.4e-07 sb=4.1e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=101380 $Y=12650 $D=28
M4259 VSS 150 4215 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.74256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=8810 $Y=46850 $D=28
M4260 4215 150 VSS VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8e-07 sb=1.26256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=9290 $Y=46850 $D=28
M4261 VSS 150 4215 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8049e-13 as=1.404e-13 pd=1.28323e-06 ps=1.14e-06 nrd=0.296664 nrs=0.230769 sa=1.28e-06 sb=7.82564e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=9770 $Y=46850 $D=28
M4262 4213 150 VSS VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.008e-13 as=1.85118e-13 pd=2.24e-06 ps=1.31613e-06 nrd=0.31375 nrs=0.289247 sa=1.7275e-06 sb=2.51e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=10330 $Y=46790 $D=28
M4263 4216 4213 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.15431e-13 pd=1.12e-06 ps=2.06077e-06 nrd=0.236842 nrs=0.372976 sa=2.81053e-07 sb=1.96947e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=11190 $Y=46830 $D=28
M4264 VSS 4213 4216 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76764e-13 as=1.368e-13 pd=1.27236e-06 ps=1.12e-06 nrd=0.306032 nrs=0.236842 sa=7.61053e-07 sb=1.95684e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=11670 $Y=46830 $D=28
M4265 4216 4213 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.72112e-13 pd=1.1e-06 ps=1.23888e-06 nrd=0.243243 nrs=0.314303 sa=1.31892e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=12230 $Y=46830 $D=28
M4266 4217 53 4216 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81e-13 as=1.332e-13 pd=1.31e-06 ps=1.1e-06 nrd=0.330533 nrs=0.243243 sa=1.79892e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=12710 $Y=46830 $D=28
M4267 4216 53 4217 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.81e-13 pd=1.1e-06 ps=1.31e-06 nrd=0.243243 nrs=0.330533 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=13270 $Y=46830 $D=28
M4268 4217 53 4216 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=13750 $Y=46830 $D=28
M4269 4215 4214 4217 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=14230 $Y=46830 $D=28
M4270 4217 4214 4215 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=14710 $Y=46830 $D=28
M4271 4215 4214 4217 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=15190 $Y=46830 $D=28
M4272 4218 53 4215 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.81838e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=15670 $Y=46830 $D=28
M4273 4215 53 4218 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.63676e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=16150 $Y=46830 $D=28
M4274 4218 53 4215 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=1.332e-13 pd=1.66e-06 ps=1.1e-06 nrd=0.514244 nrs=0.243243 sa=2e-06 sb=1.45514e-06 sd=0 panw1=0 panw2=0 panw3=6e-16 panw4=3e-15 panw5=3e-15 panw6=6.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=16630 $Y=46830 $D=28
M4275 4216 4214 4218 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.816e-13 pd=1.1e-06 ps=1.66e-06 nrd=0.243243 nrs=0.514244 sa=1.39459e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=17390 $Y=46550 $D=28
M4276 4218 4214 4216 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.09e-13 as=1.332e-13 pd=1.51e-06 ps=1.1e-06 nrd=0.381665 nrs=0.243243 sa=1.57622e-06 sb=8.8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=17870 $Y=46550 $D=28
M4277 4216 4214 4218 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=2.09e-13 pd=2.12e-06 ps=1.51e-06 nrd=0.432432 nrs=0.381665 sa=1.78811e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=18430 $Y=46550 $D=28
M4278 VSS 53 4214 VSS lpnfet w=1.07e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.93789e-13 as=3.424e-13 pd=1.76352e-06 ps=2.78e-06 nrd=0.169263 nrs=0.299065 sa=3.2e-07 sb=1.12037e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=19470 $Y=46540 $D=28
M4279 4214 53 VSS VSS lpnfet w=8.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.01576e-13 as=1.467e-13 pd=1.59826e-06 ps=1.335e-06 nrd=0.307233 nrs=0.223594 sa=7.6e-07 sb=1.19111e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=19910 $Y=46540 $D=28
M4280 VSS 53 4214 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55405e-13 as=1.69224e-13 pd=1.15268e-06 ps=1.34174e-06 nrd=0.336083 nrs=0.365969 sa=9.05294e-07 sb=1.87059e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=20430 $Y=46930 $D=28
M4281 4214 53 VSS VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30552e-13 as=1.55405e-13 pd=1.42476e-06 ps=1.15268e-06 nrd=0.498599 nrs=0.336083 sa=1.46529e-06 sb=1.44235e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=20990 $Y=46930 $D=28
M4282 4219 4217 4214 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48449e-13 as=1.96648e-13 pd=1.07378e-06 ps=1.21524e-06 nrd=0.441286 nrs=0.584565 sa=1.89517e-06 sb=8.34483e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=21750 $Y=46930 $D=28
M4283 4214 4217 4219 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.616e-13 as=2.30351e-13 pd=2.44e-06 ps=1.66622e-06 nrd=0.322963 nrs=0.284384 sa=1.41689e-06 sb=2.90667e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=22310 $Y=46610 $D=28
M4284 4219 4218 4221 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.342e-13 pd=1.12e-06 ps=2.16e-06 nrd=0.236842 nrs=0.405471 sa=3.08158e-07 sb=1.45882e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=23280 $Y=46710 $D=28
M4285 4221 4218 4219 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.52152e-13 as=1.368e-13 pd=1.3072e-06 ps=1.12e-06 nrd=0.263421 nrs=0.236842 sa=7.88158e-07 sb=9.78816e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=23760 $Y=46710 $D=28
M4286 4222 4217 4221 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.48148e-13 pd=1.1e-06 ps=1.2728e-06 nrd=0.243243 nrs=0.270541 sa=1.05027e-06 sb=7.27568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=24240 $Y=46540 $D=28
M4287 4221 4217 4222 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=1.332e-13 pd=2.8e-06 ps=1.1e-06 nrd=0.487947 nrs=0.243243 sa=1.53027e-06 sb=2.47568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=24720 $Y=46540 $D=28
M4288 4222 4218 4220 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.132e-13 pd=1.06e-06 ps=2.46e-06 nrd=0.257143 nrs=0.435102 sa=2.36571e-07 sb=1.79543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=25580 $Y=46710 $D=28
M4289 4220 4218 4222 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.16571e-07 sb=1.31543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=26060 $Y=46710 $D=28
M4290 VSS 4221 4220 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87877e-13 as=1.26e-13 pd=1.39136e-06 ps=1.06e-06 nrd=0.383422 nrs=0.257143 sa=1.19657e-06 sb=8.35429e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=26540 $Y=46710 $D=28
M4291 4220 4221 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.71773e-13 pd=1.92e-06 ps=1.2721e-06 nrd=0.5 nrs=0.419367 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=27100 $Y=46710 $D=28
M4292 VSS 94 4221 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=28040 $Y=46690 $D=28
M4293 4221 94 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=28520 $Y=46690 $D=28
M4294 44 4219 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=2.912e-13 pd=1.27e-06 ps=2.46e-06 nrd=0.197802 nrs=0.351648 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=29560 $Y=46690 $D=28
M4295 VSS 4219 44 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=1.638e-13 pd=1.27e-06 ps=1.27e-06 nrd=0.197802 nrs=0.197802 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=30040 $Y=46690 $D=28
M4296 21 4222 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=1.638e-13 pd=1.31e-06 ps=1.27e-06 nrd=0.21978 nrs=0.197802 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=30520 $Y=46690 $D=28
M4297 VSS 4222 21 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.912e-13 as=1.82e-13 pd=2.46e-06 ps=1.31e-06 nrd=0.351648 nrs=0.21978 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=31040 $Y=46690 $D=28
M4298 VSS 103 4225 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.74256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=28010 $Y=39650 $D=28
M4299 4225 103 VSS VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8e-07 sb=1.26256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=28490 $Y=39650 $D=28
M4300 VSS 103 4225 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8049e-13 as=1.404e-13 pd=1.28323e-06 ps=1.14e-06 nrd=0.296664 nrs=0.230769 sa=1.28e-06 sb=7.82564e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=28970 $Y=39650 $D=28
M4301 4223 103 VSS VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.008e-13 as=1.85118e-13 pd=2.24e-06 ps=1.31613e-06 nrd=0.31375 nrs=0.289247 sa=1.7275e-06 sb=2.51e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=29530 $Y=39590 $D=28
M4302 4226 4223 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.15431e-13 pd=1.12e-06 ps=2.06077e-06 nrd=0.236842 nrs=0.372976 sa=2.81053e-07 sb=1.96947e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=30390 $Y=39630 $D=28
M4303 VSS 4223 4226 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76764e-13 as=1.368e-13 pd=1.27236e-06 ps=1.12e-06 nrd=0.306032 nrs=0.236842 sa=7.61053e-07 sb=1.95684e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=30870 $Y=39630 $D=28
M4304 4226 4223 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.72112e-13 pd=1.1e-06 ps=1.23888e-06 nrd=0.243243 nrs=0.314303 sa=1.31892e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=31430 $Y=39630 $D=28
M4305 4227 194 4226 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81e-13 as=1.332e-13 pd=1.31e-06 ps=1.1e-06 nrd=0.330533 nrs=0.243243 sa=1.79892e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=31910 $Y=39630 $D=28
M4306 4226 194 4227 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.81e-13 pd=1.1e-06 ps=1.31e-06 nrd=0.243243 nrs=0.330533 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=32470 $Y=39630 $D=28
M4307 4227 194 4226 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=32950 $Y=39630 $D=28
M4308 4225 4224 4227 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=33430 $Y=39630 $D=28
M4309 4227 4224 4225 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=33910 $Y=39630 $D=28
M4310 4225 4224 4227 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=34390 $Y=39630 $D=28
M4311 4228 194 4225 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.81838e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=34870 $Y=39630 $D=28
M4312 4225 194 4228 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.63676e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=35350 $Y=39630 $D=28
M4313 4228 194 4225 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=1.332e-13 pd=1.66e-06 ps=1.1e-06 nrd=0.514244 nrs=0.243243 sa=2e-06 sb=1.45514e-06 sd=0 panw1=0 panw2=0 panw3=6e-16 panw4=3e-15 panw5=3e-15 panw6=6.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=35830 $Y=39630 $D=28
M4314 4226 4224 4228 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.816e-13 pd=1.1e-06 ps=1.66e-06 nrd=0.243243 nrs=0.514244 sa=1.39459e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=36590 $Y=39350 $D=28
M4315 4228 4224 4226 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.09e-13 as=1.332e-13 pd=1.51e-06 ps=1.1e-06 nrd=0.381665 nrs=0.243243 sa=1.57622e-06 sb=8.8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=37070 $Y=39350 $D=28
M4316 4226 4224 4228 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=2.09e-13 pd=2.12e-06 ps=1.51e-06 nrd=0.432432 nrs=0.381665 sa=1.78811e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=37630 $Y=39350 $D=28
M4317 VSS 194 4224 VSS lpnfet w=1.07e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.93789e-13 as=3.424e-13 pd=1.76352e-06 ps=2.78e-06 nrd=0.169263 nrs=0.299065 sa=3.2e-07 sb=1.12037e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=38670 $Y=39340 $D=28
M4318 4224 194 VSS VSS lpnfet w=8.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.01576e-13 as=1.467e-13 pd=1.59826e-06 ps=1.335e-06 nrd=0.307233 nrs=0.223594 sa=7.6e-07 sb=1.19111e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=39110 $Y=39340 $D=28
M4319 VSS 194 4224 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55405e-13 as=1.69224e-13 pd=1.15268e-06 ps=1.34174e-06 nrd=0.336083 nrs=0.365969 sa=9.05294e-07 sb=1.87059e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=39630 $Y=39730 $D=28
M4320 4224 194 VSS VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30552e-13 as=1.55405e-13 pd=1.42476e-06 ps=1.15268e-06 nrd=0.498599 nrs=0.336083 sa=1.46529e-06 sb=1.44235e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=40190 $Y=39730 $D=28
M4321 4229 4227 4224 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48449e-13 as=1.96648e-13 pd=1.07378e-06 ps=1.21524e-06 nrd=0.441286 nrs=0.584565 sa=1.89517e-06 sb=8.34483e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=40950 $Y=39730 $D=28
M4322 4224 4227 4229 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.616e-13 as=2.30351e-13 pd=2.44e-06 ps=1.66622e-06 nrd=0.322963 nrs=0.284384 sa=1.41689e-06 sb=2.90667e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=41510 $Y=39410 $D=28
M4323 4229 4228 4231 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.342e-13 pd=1.12e-06 ps=2.16e-06 nrd=0.236842 nrs=0.405471 sa=3.08158e-07 sb=1.45882e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=42480 $Y=39510 $D=28
M4324 4231 4228 4229 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.52152e-13 as=1.368e-13 pd=1.3072e-06 ps=1.12e-06 nrd=0.263421 nrs=0.236842 sa=7.88158e-07 sb=9.78816e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=42960 $Y=39510 $D=28
M4325 4232 4227 4231 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.48148e-13 pd=1.1e-06 ps=1.2728e-06 nrd=0.243243 nrs=0.270541 sa=1.05027e-06 sb=7.27568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=43440 $Y=39340 $D=28
M4326 4231 4227 4232 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=1.332e-13 pd=2.8e-06 ps=1.1e-06 nrd=0.487947 nrs=0.243243 sa=1.53027e-06 sb=2.47568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=43920 $Y=39340 $D=28
M4327 4232 4228 4230 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.132e-13 pd=1.06e-06 ps=2.46e-06 nrd=0.257143 nrs=0.435102 sa=2.36571e-07 sb=1.79543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=44780 $Y=39510 $D=28
M4328 4230 4228 4232 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.16571e-07 sb=1.31543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=45260 $Y=39510 $D=28
M4329 VSS 4231 4230 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87877e-13 as=1.26e-13 pd=1.39136e-06 ps=1.06e-06 nrd=0.383422 nrs=0.257143 sa=1.19657e-06 sb=8.35429e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=45740 $Y=39510 $D=28
M4330 4230 4231 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.71773e-13 pd=1.92e-06 ps=1.2721e-06 nrd=0.5 nrs=0.419367 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=46300 $Y=39510 $D=28
M4331 VSS 178 4231 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=47240 $Y=39490 $D=28
M4332 4231 178 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=47720 $Y=39490 $D=28
M4333 120 4229 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=2.912e-13 pd=1.27e-06 ps=2.46e-06 nrd=0.197802 nrs=0.351648 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=48760 $Y=39490 $D=28
M4334 VSS 4229 120 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=1.638e-13 pd=1.27e-06 ps=1.27e-06 nrd=0.197802 nrs=0.197802 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=49240 $Y=39490 $D=28
M4335 94 4232 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=1.638e-13 pd=1.31e-06 ps=1.27e-06 nrd=0.21978 nrs=0.197802 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=49720 $Y=39490 $D=28
M4336 VSS 4232 94 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.912e-13 as=1.82e-13 pd=2.46e-06 ps=1.31e-06 nrd=0.351648 nrs=0.21978 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=50240 $Y=39490 $D=28
M4337 VSS 253 4235 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.74256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=54010 $Y=68450 $D=28
M4338 4235 253 VSS VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8e-07 sb=1.26256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=54490 $Y=68450 $D=28
M4339 VSS 253 4235 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8049e-13 as=1.404e-13 pd=1.28323e-06 ps=1.14e-06 nrd=0.296664 nrs=0.230769 sa=1.28e-06 sb=7.82564e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=54970 $Y=68450 $D=28
M4340 4233 253 VSS VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.008e-13 as=1.85118e-13 pd=2.24e-06 ps=1.31613e-06 nrd=0.31375 nrs=0.289247 sa=1.7275e-06 sb=2.51e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=55530 $Y=68390 $D=28
M4341 4236 4233 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.15431e-13 pd=1.12e-06 ps=2.06077e-06 nrd=0.236842 nrs=0.372976 sa=2.81053e-07 sb=1.96947e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=56390 $Y=68430 $D=28
M4342 VSS 4233 4236 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76764e-13 as=1.368e-13 pd=1.27236e-06 ps=1.12e-06 nrd=0.306032 nrs=0.236842 sa=7.61053e-07 sb=1.95684e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=56870 $Y=68430 $D=28
M4343 4236 4233 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.72112e-13 pd=1.1e-06 ps=1.23888e-06 nrd=0.243243 nrs=0.314303 sa=1.31892e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=57430 $Y=68430 $D=28
M4344 4237 276 4236 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81e-13 as=1.332e-13 pd=1.31e-06 ps=1.1e-06 nrd=0.330533 nrs=0.243243 sa=1.79892e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=57910 $Y=68430 $D=28
M4345 4236 276 4237 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.81e-13 pd=1.1e-06 ps=1.31e-06 nrd=0.243243 nrs=0.330533 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=58470 $Y=68430 $D=28
M4346 4237 276 4236 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=58950 $Y=68430 $D=28
M4347 4235 4234 4237 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=59430 $Y=68430 $D=28
M4348 4237 4234 4235 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=59910 $Y=68430 $D=28
M4349 4235 4234 4237 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=60390 $Y=68430 $D=28
M4350 4238 276 4235 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.81838e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=60870 $Y=68430 $D=28
M4351 4235 276 4238 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.63676e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=61350 $Y=68430 $D=28
M4352 4238 276 4235 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=1.332e-13 pd=1.66e-06 ps=1.1e-06 nrd=0.514244 nrs=0.243243 sa=2e-06 sb=1.45514e-06 sd=0 panw1=0 panw2=0 panw3=6e-16 panw4=3e-15 panw5=3e-15 panw6=6.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=61830 $Y=68430 $D=28
M4353 4236 4234 4238 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.816e-13 pd=1.1e-06 ps=1.66e-06 nrd=0.243243 nrs=0.514244 sa=1.39459e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=62590 $Y=68150 $D=28
M4354 4238 4234 4236 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.09e-13 as=1.332e-13 pd=1.51e-06 ps=1.1e-06 nrd=0.381665 nrs=0.243243 sa=1.57622e-06 sb=8.8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=63070 $Y=68150 $D=28
M4355 4236 4234 4238 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=2.09e-13 pd=2.12e-06 ps=1.51e-06 nrd=0.432432 nrs=0.381665 sa=1.78811e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=63630 $Y=68150 $D=28
M4356 VSS 276 4234 VSS lpnfet w=1.07e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.93789e-13 as=3.424e-13 pd=1.76352e-06 ps=2.78e-06 nrd=0.169263 nrs=0.299065 sa=3.2e-07 sb=1.12037e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=64670 $Y=68140 $D=28
M4357 4234 276 VSS VSS lpnfet w=8.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.01576e-13 as=1.467e-13 pd=1.59826e-06 ps=1.335e-06 nrd=0.307233 nrs=0.223594 sa=7.6e-07 sb=1.19111e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=65110 $Y=68140 $D=28
M4358 VSS 276 4234 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55405e-13 as=1.69224e-13 pd=1.15268e-06 ps=1.34174e-06 nrd=0.336083 nrs=0.365969 sa=9.05294e-07 sb=1.87059e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=65630 $Y=68530 $D=28
M4359 4234 276 VSS VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30552e-13 as=1.55405e-13 pd=1.42476e-06 ps=1.15268e-06 nrd=0.498599 nrs=0.336083 sa=1.46529e-06 sb=1.44235e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=66190 $Y=68530 $D=28
M4360 4239 4237 4234 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48449e-13 as=1.96648e-13 pd=1.07378e-06 ps=1.21524e-06 nrd=0.441286 nrs=0.584565 sa=1.89517e-06 sb=8.34483e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=66950 $Y=68530 $D=28
M4361 4234 4237 4239 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.616e-13 as=2.30351e-13 pd=2.44e-06 ps=1.66622e-06 nrd=0.322963 nrs=0.284384 sa=1.41689e-06 sb=2.90667e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=67510 $Y=68210 $D=28
M4362 4239 4238 4241 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.342e-13 pd=1.12e-06 ps=2.16e-06 nrd=0.236842 nrs=0.405471 sa=3.08158e-07 sb=1.45882e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=68480 $Y=68310 $D=28
M4363 4241 4238 4239 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.52152e-13 as=1.368e-13 pd=1.3072e-06 ps=1.12e-06 nrd=0.263421 nrs=0.236842 sa=7.88158e-07 sb=9.78816e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=68960 $Y=68310 $D=28
M4364 4242 4237 4241 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.48148e-13 pd=1.1e-06 ps=1.2728e-06 nrd=0.243243 nrs=0.270541 sa=1.05027e-06 sb=7.27568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=69440 $Y=68140 $D=28
M4365 4241 4237 4242 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=1.332e-13 pd=2.8e-06 ps=1.1e-06 nrd=0.487947 nrs=0.243243 sa=1.53027e-06 sb=2.47568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=69920 $Y=68140 $D=28
M4366 4242 4238 4240 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.132e-13 pd=1.06e-06 ps=2.46e-06 nrd=0.257143 nrs=0.435102 sa=2.36571e-07 sb=1.79543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=70780 $Y=68310 $D=28
M4367 4240 4238 4242 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.16571e-07 sb=1.31543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=71260 $Y=68310 $D=28
M4368 VSS 4241 4240 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87877e-13 as=1.26e-13 pd=1.39136e-06 ps=1.06e-06 nrd=0.383422 nrs=0.257143 sa=1.19657e-06 sb=8.35429e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=71740 $Y=68310 $D=28
M4369 4240 4241 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.71773e-13 pd=1.92e-06 ps=1.2721e-06 nrd=0.5 nrs=0.419367 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=72300 $Y=68310 $D=28
M4370 VSS 275 4241 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=73240 $Y=68290 $D=28
M4371 4241 275 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=8e-15 $X=73720 $Y=68290 $D=28
M4372 309 4239 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=2.912e-13 pd=1.27e-06 ps=2.46e-06 nrd=0.197802 nrs=0.351648 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=1.08e-14 $X=74760 $Y=68290 $D=28
M4373 VSS 4239 309 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=1.638e-13 pd=1.27e-06 ps=1.27e-06 nrd=0.197802 nrs=0.197802 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=1.08e-14 $X=75240 $Y=68290 $D=28
M4374 289 4242 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=1.638e-13 pd=1.31e-06 ps=1.27e-06 nrd=0.21978 nrs=0.197802 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=6.3e-15 $X=75720 $Y=68290 $D=28
M4375 VSS 4242 289 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.912e-13 as=1.82e-13 pd=2.46e-06 ps=1.31e-06 nrd=0.351648 nrs=0.21978 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=76240 $Y=68290 $D=28
M4376 VSS 234 4245 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.74256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=63610 $Y=54050 $D=28
M4377 4245 234 VSS VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8e-07 sb=1.26256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=64090 $Y=54050 $D=28
M4378 VSS 234 4245 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8049e-13 as=1.404e-13 pd=1.28323e-06 ps=1.14e-06 nrd=0.296664 nrs=0.230769 sa=1.28e-06 sb=7.82564e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=64570 $Y=54050 $D=28
M4379 4243 234 VSS VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.008e-13 as=1.85118e-13 pd=2.24e-06 ps=1.31613e-06 nrd=0.31375 nrs=0.289247 sa=1.7275e-06 sb=2.51e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=65130 $Y=53990 $D=28
M4380 4246 4243 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.15431e-13 pd=1.12e-06 ps=2.06077e-06 nrd=0.236842 nrs=0.372976 sa=2.81053e-07 sb=1.96947e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=65990 $Y=54030 $D=28
M4381 VSS 4243 4246 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76764e-13 as=1.368e-13 pd=1.27236e-06 ps=1.12e-06 nrd=0.306032 nrs=0.236842 sa=7.61053e-07 sb=1.95684e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=66470 $Y=54030 $D=28
M4382 4246 4243 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.72112e-13 pd=1.1e-06 ps=1.23888e-06 nrd=0.243243 nrs=0.314303 sa=1.31892e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=67030 $Y=54030 $D=28
M4383 4247 824 4246 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81e-13 as=1.332e-13 pd=1.31e-06 ps=1.1e-06 nrd=0.330533 nrs=0.243243 sa=1.79892e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=67510 $Y=54030 $D=28
M4384 4246 824 4247 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.81e-13 pd=1.1e-06 ps=1.31e-06 nrd=0.243243 nrs=0.330533 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=68070 $Y=54030 $D=28
M4385 4247 824 4246 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=68550 $Y=54030 $D=28
M4386 4245 4244 4247 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=69030 $Y=54030 $D=28
M4387 4247 4244 4245 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=69510 $Y=54030 $D=28
M4388 4245 4244 4247 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=69990 $Y=54030 $D=28
M4389 4248 824 4245 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.81838e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=70470 $Y=54030 $D=28
M4390 4245 824 4248 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.63676e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=70950 $Y=54030 $D=28
M4391 4248 824 4245 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=1.332e-13 pd=1.66e-06 ps=1.1e-06 nrd=0.514244 nrs=0.243243 sa=2e-06 sb=1.45514e-06 sd=0 panw1=0 panw2=0 panw3=6e-16 panw4=3e-15 panw5=3e-15 panw6=6.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=71430 $Y=54030 $D=28
M4392 4246 4244 4248 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.816e-13 pd=1.1e-06 ps=1.66e-06 nrd=0.243243 nrs=0.514244 sa=1.39459e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=72190 $Y=53750 $D=28
M4393 4248 4244 4246 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.09e-13 as=1.332e-13 pd=1.51e-06 ps=1.1e-06 nrd=0.381665 nrs=0.243243 sa=1.57622e-06 sb=8.8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=72670 $Y=53750 $D=28
M4394 4246 4244 4248 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=2.09e-13 pd=2.12e-06 ps=1.51e-06 nrd=0.432432 nrs=0.381665 sa=1.78811e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=73230 $Y=53750 $D=28
M4395 VSS 824 4244 VSS lpnfet w=1.07e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.93789e-13 as=3.424e-13 pd=1.76352e-06 ps=2.78e-06 nrd=0.169263 nrs=0.299065 sa=3.2e-07 sb=1.12037e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=74270 $Y=53740 $D=28
M4396 4244 824 VSS VSS lpnfet w=8.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.01576e-13 as=1.467e-13 pd=1.59826e-06 ps=1.335e-06 nrd=0.307233 nrs=0.223594 sa=7.6e-07 sb=1.19111e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=74710 $Y=53740 $D=28
M4397 VSS 824 4244 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55405e-13 as=1.69224e-13 pd=1.15268e-06 ps=1.34174e-06 nrd=0.336083 nrs=0.365969 sa=9.05294e-07 sb=1.87059e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=75230 $Y=54130 $D=28
M4398 4244 824 VSS VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30552e-13 as=1.55405e-13 pd=1.42476e-06 ps=1.15268e-06 nrd=0.498599 nrs=0.336083 sa=1.46529e-06 sb=1.44235e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=75790 $Y=54130 $D=28
M4399 4249 4247 4244 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48449e-13 as=1.96648e-13 pd=1.07378e-06 ps=1.21524e-06 nrd=0.441286 nrs=0.584565 sa=1.89517e-06 sb=8.34483e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=76550 $Y=54130 $D=28
M4400 4244 4247 4249 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.616e-13 as=2.30351e-13 pd=2.44e-06 ps=1.66622e-06 nrd=0.322963 nrs=0.284384 sa=1.41689e-06 sb=2.90667e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=77110 $Y=53810 $D=28
M4401 4249 4248 4251 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.342e-13 pd=1.12e-06 ps=2.16e-06 nrd=0.236842 nrs=0.405471 sa=3.08158e-07 sb=1.45882e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=78080 $Y=53910 $D=28
M4402 4251 4248 4249 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.52152e-13 as=1.368e-13 pd=1.3072e-06 ps=1.12e-06 nrd=0.263421 nrs=0.236842 sa=7.88158e-07 sb=9.78816e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=78560 $Y=53910 $D=28
M4403 4252 4247 4251 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.48148e-13 pd=1.1e-06 ps=1.2728e-06 nrd=0.243243 nrs=0.270541 sa=1.05027e-06 sb=7.27568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=79040 $Y=53740 $D=28
M4404 4251 4247 4252 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=1.332e-13 pd=2.8e-06 ps=1.1e-06 nrd=0.487947 nrs=0.243243 sa=1.53027e-06 sb=2.47568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=79520 $Y=53740 $D=28
M4405 4252 4248 4250 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.132e-13 pd=1.06e-06 ps=2.46e-06 nrd=0.257143 nrs=0.435102 sa=2.36571e-07 sb=1.79543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=80380 $Y=53910 $D=28
M4406 4250 4248 4252 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.16571e-07 sb=1.31543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=80860 $Y=53910 $D=28
M4407 VSS 4251 4250 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87877e-13 as=1.26e-13 pd=1.39136e-06 ps=1.06e-06 nrd=0.383422 nrs=0.257143 sa=1.19657e-06 sb=8.35429e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=81340 $Y=53910 $D=28
M4408 4250 4251 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.71773e-13 pd=1.92e-06 ps=1.2721e-06 nrd=0.5 nrs=0.419367 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=81900 $Y=53910 $D=28
M4409 VSS 288 4251 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=82840 $Y=53890 $D=28
M4410 4251 288 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=83320 $Y=53890 $D=28
M4411 312 4249 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=2.912e-13 pd=1.27e-06 ps=2.46e-06 nrd=0.197802 nrs=0.351648 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=84360 $Y=53890 $D=28
M4412 VSS 4249 312 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=1.638e-13 pd=1.27e-06 ps=1.27e-06 nrd=0.197802 nrs=0.197802 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=84840 $Y=53890 $D=28
M4413 272 4252 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=1.638e-13 pd=1.31e-06 ps=1.27e-06 nrd=0.21978 nrs=0.197802 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=85320 $Y=53890 $D=28
M4414 VSS 4252 272 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.912e-13 as=1.82e-13 pd=2.46e-06 ps=1.31e-06 nrd=0.351648 nrs=0.21978 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=85840 $Y=53890 $D=28
M4415 VSS 312 4255 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.74256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=72010 $Y=69970 $D=28
M4416 4255 312 VSS VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8e-07 sb=1.26256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=72490 $Y=69970 $D=28
M4417 VSS 312 4255 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8049e-13 as=1.404e-13 pd=1.28323e-06 ps=1.14e-06 nrd=0.296664 nrs=0.230769 sa=1.28e-06 sb=7.82564e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=72970 $Y=69970 $D=28
M4418 4253 312 VSS VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.008e-13 as=1.85118e-13 pd=2.24e-06 ps=1.31613e-06 nrd=0.31375 nrs=0.289247 sa=1.7275e-06 sb=2.51e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=73530 $Y=70010 $D=28
M4419 4256 4253 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.15431e-13 pd=1.12e-06 ps=2.06077e-06 nrd=0.236842 nrs=0.372976 sa=2.81053e-07 sb=1.96947e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=74390 $Y=70010 $D=28
M4420 VSS 4253 4256 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76764e-13 as=1.368e-13 pd=1.27236e-06 ps=1.12e-06 nrd=0.306032 nrs=0.236842 sa=7.61053e-07 sb=1.95684e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=74870 $Y=70010 $D=28
M4421 4256 4253 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.72112e-13 pd=1.1e-06 ps=1.23888e-06 nrd=0.243243 nrs=0.314303 sa=1.31892e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=75430 $Y=70030 $D=28
M4422 4257 309 4256 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81e-13 as=1.332e-13 pd=1.31e-06 ps=1.1e-06 nrd=0.330533 nrs=0.243243 sa=1.79892e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=75910 $Y=70030 $D=28
M4423 4256 309 4257 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.81e-13 pd=1.1e-06 ps=1.31e-06 nrd=0.243243 nrs=0.330533 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=76470 $Y=70030 $D=28
M4424 4257 309 4256 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=76950 $Y=70030 $D=28
M4425 4255 4254 4257 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=77430 $Y=70030 $D=28
M4426 4257 4254 4255 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=77910 $Y=70030 $D=28
M4427 4255 4254 4257 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=78390 $Y=70030 $D=28
M4428 4258 309 4255 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.81838e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=1.8e-15 $X=78870 $Y=70030 $D=28
M4429 4255 309 4258 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.63676e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=7.2e-15 $X=79350 $Y=70030 $D=28
M4430 4258 309 4255 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=1.332e-13 pd=1.66e-06 ps=1.1e-06 nrd=0.514244 nrs=0.243243 sa=2e-06 sb=1.45514e-06 sd=0 panw1=0 panw2=0 panw3=6e-16 panw4=3e-15 panw5=3e-15 panw6=6.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=7.2e-15 $X=79830 $Y=70030 $D=28
M4431 4256 4254 4258 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.816e-13 pd=1.1e-06 ps=1.66e-06 nrd=0.243243 nrs=0.514244 sa=1.39459e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=80590 $Y=70310 $D=28
M4432 4258 4254 4256 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.09e-13 as=1.332e-13 pd=1.51e-06 ps=1.1e-06 nrd=0.381665 nrs=0.243243 sa=1.57622e-06 sb=8.8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=81070 $Y=70310 $D=28
M4433 4256 4254 4258 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=2.09e-13 pd=2.12e-06 ps=1.51e-06 nrd=0.432432 nrs=0.381665 sa=1.78811e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=81630 $Y=70310 $D=28
M4434 VSS 309 4254 VSS lpnfet w=1.07e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.93789e-13 as=3.424e-13 pd=1.76352e-06 ps=2.78e-06 nrd=0.169263 nrs=0.299065 sa=3.2e-07 sb=1.12037e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=1.2e-15 $X=82670 $Y=69990 $D=28
M4435 4254 309 VSS VSS lpnfet w=8.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.01576e-13 as=1.467e-13 pd=1.59826e-06 ps=1.335e-06 nrd=0.307233 nrs=0.223594 sa=7.6e-07 sb=1.19111e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=83110 $Y=70250 $D=28
M4436 VSS 309 4254 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55405e-13 as=1.69224e-13 pd=1.15268e-06 ps=1.34174e-06 nrd=0.336083 nrs=0.365969 sa=9.05294e-07 sb=1.87059e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=6e-15 $X=83630 $Y=69990 $D=28
M4437 4254 309 VSS VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30552e-13 as=1.55405e-13 pd=1.42476e-06 ps=1.15268e-06 nrd=0.498599 nrs=0.336083 sa=1.46529e-06 sb=1.44235e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=6e-15 $X=84190 $Y=69990 $D=28
M4438 4259 4257 4254 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48449e-13 as=1.96648e-13 pd=1.07378e-06 ps=1.21524e-06 nrd=0.441286 nrs=0.584565 sa=1.89517e-06 sb=8.34483e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=84950 $Y=70090 $D=28
M4439 4254 4257 4259 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.616e-13 as=2.30351e-13 pd=2.44e-06 ps=1.66622e-06 nrd=0.322963 nrs=0.284384 sa=1.41689e-06 sb=2.90667e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=85510 $Y=70090 $D=28
M4440 4259 4258 4261 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.342e-13 pd=1.12e-06 ps=2.16e-06 nrd=0.236842 nrs=0.405471 sa=3.08158e-07 sb=1.45882e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=86480 $Y=70130 $D=28
M4441 4261 4258 4259 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.52152e-13 as=1.368e-13 pd=1.3072e-06 ps=1.12e-06 nrd=0.263421 nrs=0.236842 sa=7.88158e-07 sb=9.78816e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=86960 $Y=70130 $D=28
M4442 4262 4257 4261 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.48148e-13 pd=1.1e-06 ps=1.2728e-06 nrd=0.243243 nrs=0.270541 sa=1.05027e-06 sb=7.27568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=87440 $Y=70320 $D=28
M4443 4261 4257 4262 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=1.332e-13 pd=2.8e-06 ps=1.1e-06 nrd=0.487947 nrs=0.243243 sa=1.53027e-06 sb=2.47568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=87920 $Y=70320 $D=28
M4444 4262 4258 4260 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.132e-13 pd=1.06e-06 ps=2.46e-06 nrd=0.257143 nrs=0.435102 sa=2.36571e-07 sb=1.79543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=88780 $Y=70190 $D=28
M4445 4260 4258 4262 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.16571e-07 sb=1.31543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=89260 $Y=70190 $D=28
M4446 VSS 4261 4260 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87877e-13 as=1.26e-13 pd=1.39136e-06 ps=1.06e-06 nrd=0.383422 nrs=0.257143 sa=1.19657e-06 sb=8.35429e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=89740 $Y=70190 $D=28
M4447 4260 4261 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.71773e-13 pd=1.92e-06 ps=1.2721e-06 nrd=0.5 nrs=0.419367 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=90300 $Y=70250 $D=28
M4448 VSS 338 4261 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=91240 $Y=69990 $D=28
M4449 4261 338 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=91720 $Y=69990 $D=28
M4450 342 4259 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=2.912e-13 pd=1.27e-06 ps=2.46e-06 nrd=0.197802 nrs=0.351648 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=92760 $Y=70000 $D=28
M4451 VSS 4259 342 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=1.638e-13 pd=1.27e-06 ps=1.27e-06 nrd=0.197802 nrs=0.197802 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=93240 $Y=70000 $D=28
M4452 347 4262 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=1.638e-13 pd=1.31e-06 ps=1.27e-06 nrd=0.21978 nrs=0.197802 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=93720 $Y=70000 $D=28
M4453 VSS 4262 347 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.912e-13 as=1.82e-13 pd=2.46e-06 ps=1.31e-06 nrd=0.351648 nrs=0.21978 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=94240 $Y=70000 $D=28
M4454 VSS 273 4265 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.74256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=72810 $Y=61250 $D=28
M4455 4265 273 VSS VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8e-07 sb=1.26256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=73290 $Y=61250 $D=28
M4456 VSS 273 4265 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8049e-13 as=1.404e-13 pd=1.28323e-06 ps=1.14e-06 nrd=0.296664 nrs=0.230769 sa=1.28e-06 sb=7.82564e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=73770 $Y=61250 $D=28
M4457 4263 273 VSS VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.008e-13 as=1.85118e-13 pd=2.24e-06 ps=1.31613e-06 nrd=0.31375 nrs=0.289247 sa=1.7275e-06 sb=2.51e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=74330 $Y=61190 $D=28
M4458 4266 4263 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.15431e-13 pd=1.12e-06 ps=2.06077e-06 nrd=0.236842 nrs=0.372976 sa=2.81053e-07 sb=1.96947e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=75190 $Y=61230 $D=28
M4459 VSS 4263 4266 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76764e-13 as=1.368e-13 pd=1.27236e-06 ps=1.12e-06 nrd=0.306032 nrs=0.236842 sa=7.61053e-07 sb=1.95684e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=75670 $Y=61230 $D=28
M4460 4266 4263 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.72112e-13 pd=1.1e-06 ps=1.23888e-06 nrd=0.243243 nrs=0.314303 sa=1.31892e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=7.2e-15 $X=76230 $Y=61230 $D=28
M4461 4267 317 4266 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81e-13 as=1.332e-13 pd=1.31e-06 ps=1.1e-06 nrd=0.330533 nrs=0.243243 sa=1.79892e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=7.2e-15 $X=76710 $Y=61230 $D=28
M4462 4266 317 4267 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.81e-13 pd=1.1e-06 ps=1.31e-06 nrd=0.243243 nrs=0.330533 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=7.2e-15 $X=77270 $Y=61230 $D=28
M4463 4267 317 4266 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=7.2e-15 $X=77750 $Y=61230 $D=28
M4464 4265 4264 4267 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=78230 $Y=61230 $D=28
M4465 4267 4264 4265 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=78710 $Y=61230 $D=28
M4466 4265 4264 4267 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=79190 $Y=61230 $D=28
M4467 4268 317 4265 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.81838e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=79670 $Y=61230 $D=28
M4468 4265 317 4268 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.63676e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=1e-16 $X=80150 $Y=61230 $D=28
M4469 4268 317 4265 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=1.332e-13 pd=1.66e-06 ps=1.1e-06 nrd=0.514244 nrs=0.243243 sa=2e-06 sb=1.45514e-06 sd=0 panw1=0 panw2=0 panw3=6e-16 panw4=3e-15 panw5=3e-15 panw6=6.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=1.2e-15 $X=80630 $Y=61230 $D=28
M4470 4266 4264 4268 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.816e-13 pd=1.1e-06 ps=1.66e-06 nrd=0.243243 nrs=0.514244 sa=1.39459e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=81390 $Y=60950 $D=28
M4471 4268 4264 4266 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.09e-13 as=1.332e-13 pd=1.51e-06 ps=1.1e-06 nrd=0.381665 nrs=0.243243 sa=1.57622e-06 sb=8.8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=81870 $Y=60950 $D=28
M4472 4266 4264 4268 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=2.09e-13 pd=2.12e-06 ps=1.51e-06 nrd=0.432432 nrs=0.381665 sa=1.78811e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=82430 $Y=60950 $D=28
M4473 VSS 317 4264 VSS lpnfet w=1.07e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.93789e-13 as=3.424e-13 pd=1.76352e-06 ps=2.78e-06 nrd=0.169263 nrs=0.299065 sa=3.2e-07 sb=1.12037e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=83470 $Y=60940 $D=28
M4474 4264 317 VSS VSS lpnfet w=8.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.01576e-13 as=1.467e-13 pd=1.59826e-06 ps=1.335e-06 nrd=0.307233 nrs=0.223594 sa=7.6e-07 sb=1.19111e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=83910 $Y=60940 $D=28
M4475 VSS 317 4264 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55405e-13 as=1.69224e-13 pd=1.15268e-06 ps=1.34174e-06 nrd=0.336083 nrs=0.365969 sa=9.05294e-07 sb=1.87059e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=84430 $Y=61330 $D=28
M4476 4264 317 VSS VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30552e-13 as=1.55405e-13 pd=1.42476e-06 ps=1.15268e-06 nrd=0.498599 nrs=0.336083 sa=1.46529e-06 sb=1.44235e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=84990 $Y=61330 $D=28
M4477 4269 4267 4264 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48449e-13 as=1.96648e-13 pd=1.07378e-06 ps=1.21524e-06 nrd=0.441286 nrs=0.584565 sa=1.89517e-06 sb=8.34483e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=85750 $Y=61330 $D=28
M4478 4264 4267 4269 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.616e-13 as=2.30351e-13 pd=2.44e-06 ps=1.66622e-06 nrd=0.322963 nrs=0.284384 sa=1.41689e-06 sb=2.90667e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=86310 $Y=61010 $D=28
M4479 4269 4268 4271 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.342e-13 pd=1.12e-06 ps=2.16e-06 nrd=0.236842 nrs=0.405471 sa=3.08158e-07 sb=1.45882e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=87280 $Y=61110 $D=28
M4480 4271 4268 4269 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.52152e-13 as=1.368e-13 pd=1.3072e-06 ps=1.12e-06 nrd=0.263421 nrs=0.236842 sa=7.88158e-07 sb=9.78816e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=87760 $Y=61110 $D=28
M4481 4272 4267 4271 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.48148e-13 pd=1.1e-06 ps=1.2728e-06 nrd=0.243243 nrs=0.270541 sa=1.05027e-06 sb=7.27568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=88240 $Y=60940 $D=28
M4482 4271 4267 4272 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=1.332e-13 pd=2.8e-06 ps=1.1e-06 nrd=0.487947 nrs=0.243243 sa=1.53027e-06 sb=2.47568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=88720 $Y=60940 $D=28
M4483 4272 4268 4270 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.132e-13 pd=1.06e-06 ps=2.46e-06 nrd=0.257143 nrs=0.435102 sa=2.36571e-07 sb=1.79543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=89580 $Y=61110 $D=28
M4484 4270 4268 4272 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.16571e-07 sb=1.31543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=90060 $Y=61110 $D=28
M4485 VSS 4271 4270 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87877e-13 as=1.26e-13 pd=1.39136e-06 ps=1.06e-06 nrd=0.383422 nrs=0.257143 sa=1.19657e-06 sb=8.35429e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=90540 $Y=61110 $D=28
M4486 4270 4271 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.71773e-13 pd=1.92e-06 ps=1.2721e-06 nrd=0.5 nrs=0.419367 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=91100 $Y=61110 $D=28
M4487 VSS 341 4271 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=92040 $Y=61090 $D=28
M4488 4271 341 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=92520 $Y=61090 $D=28
M4489 296 4269 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=2.912e-13 pd=1.27e-06 ps=2.46e-06 nrd=0.197802 nrs=0.351648 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=93560 $Y=61090 $D=28
M4490 VSS 4269 296 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=1.638e-13 pd=1.27e-06 ps=1.27e-06 nrd=0.197802 nrs=0.197802 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=94040 $Y=61090 $D=28
M4491 829 4272 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=1.638e-13 pd=1.31e-06 ps=1.27e-06 nrd=0.21978 nrs=0.197802 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=94520 $Y=61090 $D=28
M4492 VSS 4272 829 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.912e-13 as=1.82e-13 pd=2.46e-06 ps=1.31e-06 nrd=0.351648 nrs=0.21978 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=95040 $Y=61090 $D=28
M4493 VSS 311 4275 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.74256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=74410 $Y=62770 $D=28
M4494 4275 311 VSS VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8e-07 sb=1.26256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=1.44e-14 $X=74890 $Y=62770 $D=28
M4495 VSS 311 4275 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8049e-13 as=1.404e-13 pd=1.28323e-06 ps=1.14e-06 nrd=0.296664 nrs=0.230769 sa=1.28e-06 sb=7.82564e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=1.44e-14 $X=75370 $Y=62770 $D=28
M4496 4273 311 VSS VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.008e-13 as=1.85118e-13 pd=2.24e-06 ps=1.31613e-06 nrd=0.31375 nrs=0.289247 sa=1.7275e-06 sb=2.51e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=9.6e-15 $X=75930 $Y=62810 $D=28
M4497 4276 4273 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.15431e-13 pd=1.12e-06 ps=2.06077e-06 nrd=0.236842 nrs=0.372976 sa=2.81053e-07 sb=1.96947e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=76790 $Y=62810 $D=28
M4498 VSS 4273 4276 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76764e-13 as=1.368e-13 pd=1.27236e-06 ps=1.12e-06 nrd=0.306032 nrs=0.236842 sa=7.61053e-07 sb=1.95684e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=77270 $Y=62810 $D=28
M4499 4276 4273 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.72112e-13 pd=1.1e-06 ps=1.23888e-06 nrd=0.243243 nrs=0.314303 sa=1.31892e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=77830 $Y=62830 $D=28
M4500 4277 315 4276 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81e-13 as=1.332e-13 pd=1.31e-06 ps=1.1e-06 nrd=0.330533 nrs=0.243243 sa=1.79892e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=78310 $Y=62830 $D=28
M4501 4276 315 4277 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.81e-13 pd=1.1e-06 ps=1.31e-06 nrd=0.243243 nrs=0.330533 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=1.2e-15 $X=78870 $Y=62830 $D=28
M4502 4277 315 4276 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=1.2e-15 $X=79350 $Y=62830 $D=28
M4503 4275 4274 4277 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=1.2e-15 $X=79830 $Y=62830 $D=28
M4504 4277 4274 4275 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=1.2e-15 $X=80310 $Y=62830 $D=28
M4505 4275 4274 4277 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=80790 $Y=62830 $D=28
M4506 4278 315 4275 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.81838e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=81270 $Y=62830 $D=28
M4507 4275 315 4278 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.63676e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=81750 $Y=62830 $D=28
M4508 4278 315 4275 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=1.332e-13 pd=1.66e-06 ps=1.1e-06 nrd=0.514244 nrs=0.243243 sa=2e-06 sb=1.45514e-06 sd=0 panw1=0 panw2=0 panw3=6e-16 panw4=3e-15 panw5=3e-15 panw6=6.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=82230 $Y=62830 $D=28
M4509 4276 4274 4278 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.816e-13 pd=1.1e-06 ps=1.66e-06 nrd=0.243243 nrs=0.514244 sa=1.39459e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=82990 $Y=63110 $D=28
M4510 4278 4274 4276 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.09e-13 as=1.332e-13 pd=1.51e-06 ps=1.1e-06 nrd=0.381665 nrs=0.243243 sa=1.57622e-06 sb=8.8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=83470 $Y=63110 $D=28
M4511 4276 4274 4278 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=2.09e-13 pd=2.12e-06 ps=1.51e-06 nrd=0.432432 nrs=0.381665 sa=1.78811e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=84030 $Y=63110 $D=28
M4512 VSS 315 4274 VSS lpnfet w=1.07e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.93789e-13 as=3.424e-13 pd=1.76352e-06 ps=2.78e-06 nrd=0.169263 nrs=0.299065 sa=3.2e-07 sb=1.12037e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=85070 $Y=62790 $D=28
M4513 4274 315 VSS VSS lpnfet w=8.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.01576e-13 as=1.467e-13 pd=1.59826e-06 ps=1.335e-06 nrd=0.307233 nrs=0.223594 sa=7.6e-07 sb=1.19111e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=85510 $Y=63050 $D=28
M4514 VSS 315 4274 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55405e-13 as=1.69224e-13 pd=1.15268e-06 ps=1.34174e-06 nrd=0.336083 nrs=0.365969 sa=9.05294e-07 sb=1.87059e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=86030 $Y=62790 $D=28
M4515 4274 315 VSS VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30552e-13 as=1.55405e-13 pd=1.42476e-06 ps=1.15268e-06 nrd=0.498599 nrs=0.336083 sa=1.46529e-06 sb=1.44235e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=86590 $Y=62790 $D=28
M4516 4279 4277 4274 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48449e-13 as=1.96648e-13 pd=1.07378e-06 ps=1.21524e-06 nrd=0.441286 nrs=0.584565 sa=1.89517e-06 sb=8.34483e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=87350 $Y=62890 $D=28
M4517 4274 4277 4279 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.616e-13 as=2.30351e-13 pd=2.44e-06 ps=1.66622e-06 nrd=0.322963 nrs=0.284384 sa=1.41689e-06 sb=2.90667e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=87910 $Y=62890 $D=28
M4518 4279 4278 4281 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.342e-13 pd=1.12e-06 ps=2.16e-06 nrd=0.236842 nrs=0.405471 sa=3.08158e-07 sb=1.45882e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=88880 $Y=62930 $D=28
M4519 4281 4278 4279 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.52152e-13 as=1.368e-13 pd=1.3072e-06 ps=1.12e-06 nrd=0.263421 nrs=0.236842 sa=7.88158e-07 sb=9.78816e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=89360 $Y=62930 $D=28
M4520 4282 4277 4281 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.48148e-13 pd=1.1e-06 ps=1.2728e-06 nrd=0.243243 nrs=0.270541 sa=1.05027e-06 sb=7.27568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=89840 $Y=63120 $D=28
M4521 4281 4277 4282 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=1.332e-13 pd=2.8e-06 ps=1.1e-06 nrd=0.487947 nrs=0.243243 sa=1.53027e-06 sb=2.47568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=90320 $Y=63120 $D=28
M4522 4282 4278 4280 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.132e-13 pd=1.06e-06 ps=2.46e-06 nrd=0.257143 nrs=0.435102 sa=2.36571e-07 sb=1.79543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=91180 $Y=62990 $D=28
M4523 4280 4278 4282 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.16571e-07 sb=1.31543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=91660 $Y=62990 $D=28
M4524 VSS 4281 4280 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87877e-13 as=1.26e-13 pd=1.39136e-06 ps=1.06e-06 nrd=0.383422 nrs=0.257143 sa=1.19657e-06 sb=8.35429e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=92140 $Y=62990 $D=28
M4525 4280 4281 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.71773e-13 pd=1.92e-06 ps=1.2721e-06 nrd=0.5 nrs=0.419367 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=92700 $Y=63050 $D=28
M4526 VSS 829 4281 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=93640 $Y=62790 $D=28
M4527 4281 829 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=94120 $Y=62790 $D=28
M4528 349 4279 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=2.912e-13 pd=1.27e-06 ps=2.46e-06 nrd=0.197802 nrs=0.351648 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=95160 $Y=62800 $D=28
M4529 VSS 4279 349 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=1.638e-13 pd=1.27e-06 ps=1.27e-06 nrd=0.197802 nrs=0.197802 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=95640 $Y=62800 $D=28
M4530 338 4282 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=1.638e-13 pd=1.31e-06 ps=1.27e-06 nrd=0.21978 nrs=0.197802 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=96120 $Y=62800 $D=28
M4531 VSS 4282 338 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.912e-13 as=1.82e-13 pd=2.46e-06 ps=1.31e-06 nrd=0.351648 nrs=0.21978 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=96640 $Y=62800 $D=28
M4532 VSS 296 4285 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.74256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=3.6e-15 $X=77210 $Y=68450 $D=28
M4533 4285 296 VSS VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8e-07 sb=1.26256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=3.6e-15 $X=77690 $Y=68450 $D=28
M4534 VSS 296 4285 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8049e-13 as=1.404e-13 pd=1.28323e-06 ps=1.14e-06 nrd=0.296664 nrs=0.230769 sa=1.28e-06 sb=7.82564e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=8.4e-15 $X=78170 $Y=68450 $D=28
M4535 4283 296 VSS VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.008e-13 as=1.85118e-13 pd=2.24e-06 ps=1.31613e-06 nrd=0.31375 nrs=0.289247 sa=1.7275e-06 sb=2.51e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=3.6e-15 $X=78730 $Y=68390 $D=28
M4536 4286 4283 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.15431e-13 pd=1.12e-06 ps=2.06077e-06 nrd=0.236842 nrs=0.372976 sa=2.81053e-07 sb=1.96947e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=3.6e-15 $X=79590 $Y=68430 $D=28
M4537 VSS 4283 4286 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76764e-13 as=1.368e-13 pd=1.27236e-06 ps=1.12e-06 nrd=0.306032 nrs=0.236842 sa=7.61053e-07 sb=1.95684e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=80070 $Y=68430 $D=28
M4538 4286 4283 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.72112e-13 pd=1.1e-06 ps=1.23888e-06 nrd=0.243243 nrs=0.314303 sa=1.31892e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=80630 $Y=68430 $D=28
M4539 4287 349 4286 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81e-13 as=1.332e-13 pd=1.31e-06 ps=1.1e-06 nrd=0.330533 nrs=0.243243 sa=1.79892e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=81110 $Y=68430 $D=28
M4540 4286 349 4287 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.81e-13 pd=1.1e-06 ps=1.31e-06 nrd=0.243243 nrs=0.330533 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=81670 $Y=68430 $D=28
M4541 4287 349 4286 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=82150 $Y=68430 $D=28
M4542 4285 4284 4287 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=82630 $Y=68430 $D=28
M4543 4287 4284 4285 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=83110 $Y=68430 $D=28
M4544 4285 4284 4287 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=83590 $Y=68430 $D=28
M4545 4288 349 4285 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.81838e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=84070 $Y=68430 $D=28
M4546 4285 349 4288 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.63676e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=84550 $Y=68430 $D=28
M4547 4288 349 4285 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=1.332e-13 pd=1.66e-06 ps=1.1e-06 nrd=0.514244 nrs=0.243243 sa=2e-06 sb=1.45514e-06 sd=0 panw1=0 panw2=0 panw3=6e-16 panw4=3e-15 panw5=3e-15 panw6=6.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=85030 $Y=68430 $D=28
M4548 4286 4284 4288 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.816e-13 pd=1.1e-06 ps=1.66e-06 nrd=0.243243 nrs=0.514244 sa=1.39459e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=85790 $Y=68150 $D=28
M4549 4288 4284 4286 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.09e-13 as=1.332e-13 pd=1.51e-06 ps=1.1e-06 nrd=0.381665 nrs=0.243243 sa=1.57622e-06 sb=8.8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=86270 $Y=68150 $D=28
M4550 4286 4284 4288 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=2.09e-13 pd=2.12e-06 ps=1.51e-06 nrd=0.432432 nrs=0.381665 sa=1.78811e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=86830 $Y=68150 $D=28
M4551 VSS 349 4284 VSS lpnfet w=1.07e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.93789e-13 as=3.424e-13 pd=1.76352e-06 ps=2.78e-06 nrd=0.169263 nrs=0.299065 sa=3.2e-07 sb=1.12037e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=87870 $Y=68140 $D=28
M4552 4284 349 VSS VSS lpnfet w=8.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.01576e-13 as=1.467e-13 pd=1.59826e-06 ps=1.335e-06 nrd=0.307233 nrs=0.223594 sa=7.6e-07 sb=1.19111e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=88310 $Y=68140 $D=28
M4553 VSS 349 4284 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55405e-13 as=1.69224e-13 pd=1.15268e-06 ps=1.34174e-06 nrd=0.336083 nrs=0.365969 sa=9.05294e-07 sb=1.87059e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=88830 $Y=68530 $D=28
M4554 4284 349 VSS VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30552e-13 as=1.55405e-13 pd=1.42476e-06 ps=1.15268e-06 nrd=0.498599 nrs=0.336083 sa=1.46529e-06 sb=1.44235e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=89390 $Y=68530 $D=28
M4555 4289 4287 4284 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48449e-13 as=1.96648e-13 pd=1.07378e-06 ps=1.21524e-06 nrd=0.441286 nrs=0.584565 sa=1.89517e-06 sb=8.34483e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=90150 $Y=68530 $D=28
M4556 4284 4287 4289 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.616e-13 as=2.30351e-13 pd=2.44e-06 ps=1.66622e-06 nrd=0.322963 nrs=0.284384 sa=1.41689e-06 sb=2.90667e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=90710 $Y=68210 $D=28
M4557 4289 4288 4291 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.342e-13 pd=1.12e-06 ps=2.16e-06 nrd=0.236842 nrs=0.405471 sa=3.08158e-07 sb=1.45882e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=91680 $Y=68310 $D=28
M4558 4291 4288 4289 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.52152e-13 as=1.368e-13 pd=1.3072e-06 ps=1.12e-06 nrd=0.263421 nrs=0.236842 sa=7.88158e-07 sb=9.78816e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=92160 $Y=68310 $D=28
M4559 4292 4287 4291 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.48148e-13 pd=1.1e-06 ps=1.2728e-06 nrd=0.243243 nrs=0.270541 sa=1.05027e-06 sb=7.27568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=92640 $Y=68140 $D=28
M4560 4291 4287 4292 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=1.332e-13 pd=2.8e-06 ps=1.1e-06 nrd=0.487947 nrs=0.243243 sa=1.53027e-06 sb=2.47568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=93120 $Y=68140 $D=28
M4561 4292 4288 4290 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.132e-13 pd=1.06e-06 ps=2.46e-06 nrd=0.257143 nrs=0.435102 sa=2.36571e-07 sb=1.79543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=93980 $Y=68310 $D=28
M4562 4290 4288 4292 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.16571e-07 sb=1.31543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=94460 $Y=68310 $D=28
M4563 VSS 4291 4290 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87877e-13 as=1.26e-13 pd=1.39136e-06 ps=1.06e-06 nrd=0.383422 nrs=0.257143 sa=1.19657e-06 sb=8.35429e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=94940 $Y=68310 $D=28
M4564 4290 4291 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.71773e-13 pd=1.92e-06 ps=1.2721e-06 nrd=0.5 nrs=0.419367 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=95500 $Y=68310 $D=28
M4565 VSS 831 4291 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=96440 $Y=68290 $D=28
M4566 4291 831 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=96920 $Y=68290 $D=28
M4567 401 4289 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=2.912e-13 pd=1.27e-06 ps=2.46e-06 nrd=0.197802 nrs=0.351648 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=97960 $Y=68290 $D=28
M4568 VSS 4289 401 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=1.638e-13 pd=1.27e-06 ps=1.27e-06 nrd=0.197802 nrs=0.197802 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=98440 $Y=68290 $D=28
M4569 323 4292 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=1.638e-13 pd=1.31e-06 ps=1.27e-06 nrd=0.21978 nrs=0.197802 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=98920 $Y=68290 $D=28
M4570 VSS 4292 323 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.912e-13 as=1.82e-13 pd=2.46e-06 ps=1.31e-06 nrd=0.351648 nrs=0.21978 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=99440 $Y=68290 $D=28
M4571 VSS 365 4295 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.74256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=95610 $Y=39650 $D=28
M4572 4295 365 VSS VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8e-07 sb=1.26256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=96090 $Y=39650 $D=28
M4573 VSS 365 4295 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8049e-13 as=1.404e-13 pd=1.28323e-06 ps=1.14e-06 nrd=0.296664 nrs=0.230769 sa=1.28e-06 sb=7.82564e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=96570 $Y=39650 $D=28
M4574 4293 365 VSS VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.008e-13 as=1.85118e-13 pd=2.24e-06 ps=1.31613e-06 nrd=0.31375 nrs=0.289247 sa=1.7275e-06 sb=2.51e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=97130 $Y=39590 $D=28
M4575 4296 4293 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.15431e-13 pd=1.12e-06 ps=2.06077e-06 nrd=0.236842 nrs=0.372976 sa=2.81053e-07 sb=1.96947e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=97990 $Y=39630 $D=28
M4576 VSS 4293 4296 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76764e-13 as=1.368e-13 pd=1.27236e-06 ps=1.12e-06 nrd=0.306032 nrs=0.236842 sa=7.61053e-07 sb=1.95684e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=98470 $Y=39630 $D=28
M4577 4296 4293 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.72112e-13 pd=1.1e-06 ps=1.23888e-06 nrd=0.243243 nrs=0.314303 sa=1.31892e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=99030 $Y=39630 $D=28
M4578 4297 350 4296 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81e-13 as=1.332e-13 pd=1.31e-06 ps=1.1e-06 nrd=0.330533 nrs=0.243243 sa=1.79892e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=99510 $Y=39630 $D=28
M4579 4296 350 4297 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.81e-13 pd=1.1e-06 ps=1.31e-06 nrd=0.243243 nrs=0.330533 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=100070 $Y=39630 $D=28
M4580 4297 350 4296 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=100550 $Y=39630 $D=28
M4581 4295 4294 4297 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=101030 $Y=39630 $D=28
M4582 4297 4294 4295 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=101510 $Y=39630 $D=28
M4583 4295 4294 4297 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=101990 $Y=39630 $D=28
M4584 4298 350 4295 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.81838e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=102470 $Y=39630 $D=28
M4585 4295 350 4298 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.63676e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=102950 $Y=39630 $D=28
M4586 4298 350 4295 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=1.332e-13 pd=1.66e-06 ps=1.1e-06 nrd=0.514244 nrs=0.243243 sa=2e-06 sb=1.45514e-06 sd=0 panw1=0 panw2=0 panw3=6e-16 panw4=3e-15 panw5=3e-15 panw6=6.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=103430 $Y=39630 $D=28
M4587 4296 4294 4298 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.816e-13 pd=1.1e-06 ps=1.66e-06 nrd=0.243243 nrs=0.514244 sa=1.39459e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=104190 $Y=39350 $D=28
M4588 4298 4294 4296 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.09e-13 as=1.332e-13 pd=1.51e-06 ps=1.1e-06 nrd=0.381665 nrs=0.243243 sa=1.57622e-06 sb=8.8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=104670 $Y=39350 $D=28
M4589 4296 4294 4298 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=2.09e-13 pd=2.12e-06 ps=1.51e-06 nrd=0.432432 nrs=0.381665 sa=1.78811e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=105230 $Y=39350 $D=28
M4590 VSS 350 4294 VSS lpnfet w=1.07e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.93789e-13 as=3.424e-13 pd=1.76352e-06 ps=2.78e-06 nrd=0.169263 nrs=0.299065 sa=3.2e-07 sb=1.12037e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=106270 $Y=39340 $D=28
M4591 4294 350 VSS VSS lpnfet w=8.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.01576e-13 as=1.467e-13 pd=1.59826e-06 ps=1.335e-06 nrd=0.307233 nrs=0.223594 sa=7.6e-07 sb=1.19111e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=106710 $Y=39340 $D=28
M4592 VSS 350 4294 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55405e-13 as=1.69224e-13 pd=1.15268e-06 ps=1.34174e-06 nrd=0.336083 nrs=0.365969 sa=9.05294e-07 sb=1.87059e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=107230 $Y=39730 $D=28
M4593 4294 350 VSS VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30552e-13 as=1.55405e-13 pd=1.42476e-06 ps=1.15268e-06 nrd=0.498599 nrs=0.336083 sa=1.46529e-06 sb=1.44235e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=107790 $Y=39730 $D=28
M4594 4299 4297 4294 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48449e-13 as=1.96648e-13 pd=1.07378e-06 ps=1.21524e-06 nrd=0.441286 nrs=0.584565 sa=1.89517e-06 sb=8.34483e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=108550 $Y=39730 $D=28
M4595 4294 4297 4299 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.616e-13 as=2.30351e-13 pd=2.44e-06 ps=1.66622e-06 nrd=0.322963 nrs=0.284384 sa=1.41689e-06 sb=2.90667e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=109110 $Y=39410 $D=28
M4596 4299 4298 4301 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.342e-13 pd=1.12e-06 ps=2.16e-06 nrd=0.236842 nrs=0.405471 sa=3.08158e-07 sb=1.45882e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=110080 $Y=39510 $D=28
M4597 4301 4298 4299 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.52152e-13 as=1.368e-13 pd=1.3072e-06 ps=1.12e-06 nrd=0.263421 nrs=0.236842 sa=7.88158e-07 sb=9.78816e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=110560 $Y=39510 $D=28
M4598 4302 4297 4301 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.48148e-13 pd=1.1e-06 ps=1.2728e-06 nrd=0.243243 nrs=0.270541 sa=1.05027e-06 sb=7.27568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=111040 $Y=39340 $D=28
M4599 4301 4297 4302 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=1.332e-13 pd=2.8e-06 ps=1.1e-06 nrd=0.487947 nrs=0.243243 sa=1.53027e-06 sb=2.47568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=111520 $Y=39340 $D=28
M4600 4302 4298 4300 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.132e-13 pd=1.06e-06 ps=2.46e-06 nrd=0.257143 nrs=0.435102 sa=2.36571e-07 sb=1.79543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=112380 $Y=39510 $D=28
M4601 4300 4298 4302 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.16571e-07 sb=1.31543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=112860 $Y=39510 $D=28
M4602 VSS 4301 4300 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87877e-13 as=1.26e-13 pd=1.39136e-06 ps=1.06e-06 nrd=0.383422 nrs=0.257143 sa=1.19657e-06 sb=8.35429e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=113340 $Y=39510 $D=28
M4603 4300 4301 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.71773e-13 pd=1.92e-06 ps=1.2721e-06 nrd=0.5 nrs=0.419367 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=113900 $Y=39510 $D=28
M4604 VSS 837 4301 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=114840 $Y=39490 $D=28
M4605 4301 837 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=115320 $Y=39490 $D=28
M4606 461 4299 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=2.912e-13 pd=1.27e-06 ps=2.46e-06 nrd=0.197802 nrs=0.351648 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=116360 $Y=39490 $D=28
M4607 VSS 4299 461 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=1.638e-13 pd=1.27e-06 ps=1.27e-06 nrd=0.197802 nrs=0.197802 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=116840 $Y=39490 $D=28
M4608 434 4302 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=1.638e-13 pd=1.31e-06 ps=1.27e-06 nrd=0.21978 nrs=0.197802 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=117320 $Y=39490 $D=28
M4609 VSS 4302 434 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.912e-13 as=1.82e-13 pd=2.46e-06 ps=1.31e-06 nrd=0.351648 nrs=0.21978 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=117840 $Y=39490 $D=28
M4610 VSS 382 4305 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.74256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=100410 $Y=68450 $D=28
M4611 4305 382 VSS VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8e-07 sb=1.26256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=100890 $Y=68450 $D=28
M4612 VSS 382 4305 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8049e-13 as=1.404e-13 pd=1.28323e-06 ps=1.14e-06 nrd=0.296664 nrs=0.230769 sa=1.28e-06 sb=7.82564e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=4.8e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=2.4e-15 $X=101370 $Y=68450 $D=28
M4613 4303 382 VSS VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.008e-13 as=1.85118e-13 pd=2.24e-06 ps=1.31613e-06 nrd=0.31375 nrs=0.289247 sa=1.7275e-06 sb=2.51e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=101930 $Y=68390 $D=28
M4614 4306 4303 VSS VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.15431e-13 pd=1.12e-06 ps=2.06077e-06 nrd=0.236842 nrs=0.372976 sa=2.81053e-07 sb=1.96947e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=102790 $Y=68430 $D=28
M4615 VSS 4303 4306 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.76764e-13 as=1.368e-13 pd=1.27236e-06 ps=1.12e-06 nrd=0.306032 nrs=0.236842 sa=7.61053e-07 sb=1.95684e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=103270 $Y=68430 $D=28
M4616 4306 4303 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.72112e-13 pd=1.1e-06 ps=1.23888e-06 nrd=0.243243 nrs=0.314303 sa=1.31892e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=103830 $Y=68430 $D=28
M4617 4307 434 4306 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81e-13 as=1.332e-13 pd=1.31e-06 ps=1.1e-06 nrd=0.330533 nrs=0.243243 sa=1.79892e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=104310 $Y=68430 $D=28
M4618 4306 434 4307 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.81e-13 pd=1.1e-06 ps=1.31e-06 nrd=0.243243 nrs=0.330533 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=104870 $Y=68430 $D=28
M4619 4307 434 4306 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=105350 $Y=68430 $D=28
M4620 4305 4304 4307 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=105830 $Y=68430 $D=28
M4621 4307 4304 4305 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=106310 $Y=68430 $D=28
M4622 4305 4304 4307 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=106790 $Y=68430 $D=28
M4623 4308 434 4305 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.81838e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=107270 $Y=68430 $D=28
M4624 4305 434 4308 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.332e-13 pd=1.1e-06 ps=1.1e-06 nrd=0.243243 nrs=0.243243 sa=2e-06 sb=1.63676e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=107750 $Y=68430 $D=28
M4625 4308 434 4305 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=1.332e-13 pd=1.66e-06 ps=1.1e-06 nrd=0.514244 nrs=0.243243 sa=2e-06 sb=1.45514e-06 sd=0 panw1=0 panw2=0 panw3=6e-16 panw4=3e-15 panw5=3e-15 panw6=6.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=108230 $Y=68430 $D=28
M4626 4306 4304 4308 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=2.816e-13 pd=1.1e-06 ps=1.66e-06 nrd=0.243243 nrs=0.514244 sa=1.39459e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=108990 $Y=68150 $D=28
M4627 4308 4304 4306 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.09e-13 as=1.332e-13 pd=1.51e-06 ps=1.1e-06 nrd=0.381665 nrs=0.243243 sa=1.57622e-06 sb=8.8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=109470 $Y=68150 $D=28
M4628 4306 4304 4308 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=2.09e-13 pd=2.12e-06 ps=1.51e-06 nrd=0.432432 nrs=0.381665 sa=1.78811e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6e-15 panw10=0 $X=110030 $Y=68150 $D=28
M4629 VSS 434 4304 VSS lpnfet w=1.07e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.93789e-13 as=3.424e-13 pd=1.76352e-06 ps=2.78e-06 nrd=0.169263 nrs=0.299065 sa=3.2e-07 sb=1.12037e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=111070 $Y=68140 $D=28
M4630 4304 434 VSS VSS lpnfet w=8.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.01576e-13 as=1.467e-13 pd=1.59826e-06 ps=1.335e-06 nrd=0.307233 nrs=0.223594 sa=7.6e-07 sb=1.19111e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=111510 $Y=68140 $D=28
M4631 VSS 434 4304 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55405e-13 as=1.69224e-13 pd=1.15268e-06 ps=1.34174e-06 nrd=0.336083 nrs=0.365969 sa=9.05294e-07 sb=1.87059e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=112030 $Y=68530 $D=28
M4632 4304 434 VSS VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30552e-13 as=1.55405e-13 pd=1.42476e-06 ps=1.15268e-06 nrd=0.498599 nrs=0.336083 sa=1.46529e-06 sb=1.44235e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=4.44e-14 panw10=0 $X=112590 $Y=68530 $D=28
M4633 4309 4307 4304 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48449e-13 as=1.96648e-13 pd=1.07378e-06 ps=1.21524e-06 nrd=0.441286 nrs=0.584565 sa=1.89517e-06 sb=8.34483e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.32e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=113350 $Y=68530 $D=28
M4634 4304 4307 4309 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.616e-13 as=2.30351e-13 pd=2.44e-06 ps=1.66622e-06 nrd=0.322963 nrs=0.284384 sa=1.41689e-06 sb=2.90667e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=113910 $Y=68210 $D=28
M4635 4309 4308 4311 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.368e-13 as=2.342e-13 pd=1.12e-06 ps=2.16e-06 nrd=0.236842 nrs=0.405471 sa=3.08158e-07 sb=1.45882e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=114880 $Y=68310 $D=28
M4636 4311 4308 4309 VSS lpnfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.52152e-13 as=1.368e-13 pd=1.3072e-06 ps=1.12e-06 nrd=0.263421 nrs=0.236842 sa=7.88158e-07 sb=9.78816e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=115360 $Y=68310 $D=28
M4637 4312 4307 4311 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.332e-13 as=1.48148e-13 pd=1.1e-06 ps=1.2728e-06 nrd=0.243243 nrs=0.270541 sa=1.05027e-06 sb=7.27568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=115840 $Y=68140 $D=28
M4638 4311 4307 4312 VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.672e-13 as=1.332e-13 pd=2.8e-06 ps=1.1e-06 nrd=0.487947 nrs=0.243243 sa=1.53027e-06 sb=2.47568e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=116320 $Y=68140 $D=28
M4639 4312 4308 4310 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=2.132e-13 pd=1.06e-06 ps=2.46e-06 nrd=0.257143 nrs=0.435102 sa=2.36571e-07 sb=1.79543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=117180 $Y=68310 $D=28
M4640 4310 4308 4312 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=7.16571e-07 sb=1.31543e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=117660 $Y=68310 $D=28
M4641 VSS 4311 4310 VSS lpnfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87877e-13 as=1.26e-13 pd=1.39136e-06 ps=1.06e-06 nrd=0.383422 nrs=0.257143 sa=1.19657e-06 sb=8.35429e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=118140 $Y=68310 $D=28
M4642 4310 4311 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.71773e-13 pd=1.92e-06 ps=1.2721e-06 nrd=0.5 nrs=0.419367 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=118700 $Y=68310 $D=28
M4643 VSS 381 4311 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.944e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.347826 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=119640 $Y=68290 $D=28
M4644 4311 381 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=120120 $Y=68290 $D=28
M4645 433 4309 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=2.912e-13 pd=1.27e-06 ps=2.46e-06 nrd=0.197802 nrs=0.351648 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=121160 $Y=68290 $D=28
M4646 VSS 4309 433 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=1.638e-13 pd=1.27e-06 ps=1.27e-06 nrd=0.197802 nrs=0.197802 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=121640 $Y=68290 $D=28
M4647 392 4312 VSS VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=1.638e-13 pd=1.31e-06 ps=1.27e-06 nrd=0.21978 nrs=0.197802 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=122120 $Y=68290 $D=28
M4648 VSS 4312 392 VSS lpnfet w=9.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.912e-13 as=1.82e-13 pd=2.46e-06 ps=1.31e-06 nrd=0.351648 nrs=0.21978 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=122640 $Y=68290 $D=28
M4649 VSS 35 4313 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55077e-14 as=9.6e-14 pd=5.41538e-07 ps=1.28e-06 nrd=1.14685 nrs=1.98347 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=10850 $Y=49090 $D=28
M4650 4315 13 VSS VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.41292e-13 pd=9.2e-07 ps=1.37846e-06 nrd=0.321429 nrs=0.450549 sa=5.4e-07 sb=1.96e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=11370 $Y=48750 $D=28
M4651 28 4313 4315 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.008e-13 pd=9.2e-07 ps=9.2e-07 nrd=0.321429 nrs=0.321429 sa=1.02e-06 sb=1.48e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=11850 $Y=48750 $D=28
M4652 4314 35 28 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.456e-13 as=1.008e-13 pd=1.08e-06 ps=9.2e-07 nrd=0.464286 nrs=0.321429 sa=1.5e-06 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=12330 $Y=48750 $D=28
M4653 VSS 4315 4314 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.52e-13 as=1.456e-13 pd=2.06667e-06 ps=1.08e-06 nrd=0.803571 nrs=0.464286 sa=1.95143e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=12970 $Y=48750 $D=28
M4654 VSS 19 4316 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55077e-14 as=9.6e-14 pd=5.41538e-07 ps=1.28e-06 nrd=1.14685 nrs=1.98347 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=11250 $Y=17890 $D=28
M4655 4318 15 VSS VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.41292e-13 pd=9.2e-07 ps=1.37846e-06 nrd=0.321429 nrs=0.450549 sa=5.4e-07 sb=1.96e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=11770 $Y=17890 $D=28
M4656 10 4316 4318 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.008e-13 pd=9.2e-07 ps=9.2e-07 nrd=0.321429 nrs=0.321429 sa=1.02e-06 sb=1.48e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=12250 $Y=17890 $D=28
M4657 4317 19 10 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.456e-13 as=1.008e-13 pd=1.08e-06 ps=9.2e-07 nrd=0.464286 nrs=0.321429 sa=1.5e-06 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=12730 $Y=17890 $D=28
M4658 VSS 4318 4317 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.52e-13 as=1.456e-13 pd=2.06667e-06 ps=1.08e-06 nrd=0.803571 nrs=0.464286 sa=1.95143e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=13370 $Y=17890 $D=28
M4659 VSS 802 4319 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55077e-14 as=9.6e-14 pd=5.41538e-07 ps=1.28e-06 nrd=1.14685 nrs=1.98347 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=18050 $Y=70690 $D=28
M4660 4321 64 VSS VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.41292e-13 pd=9.2e-07 ps=1.37846e-06 nrd=0.321429 nrs=0.450549 sa=5.4e-07 sb=1.96e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=18570 $Y=70350 $D=28
M4661 55 4319 4321 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.008e-13 pd=9.2e-07 ps=9.2e-07 nrd=0.321429 nrs=0.321429 sa=1.02e-06 sb=1.48e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=19050 $Y=70350 $D=28
M4662 4320 802 55 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.456e-13 as=1.008e-13 pd=1.08e-06 ps=9.2e-07 nrd=0.464286 nrs=0.321429 sa=1.5e-06 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=19530 $Y=70350 $D=28
M4663 VSS 4321 4320 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.52e-13 as=1.456e-13 pd=2.06667e-06 ps=1.08e-06 nrd=0.803571 nrs=0.464286 sa=1.95143e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=20170 $Y=70350 $D=28
M4664 VSS 101 4322 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55077e-14 as=9.6e-14 pd=5.41538e-07 ps=1.28e-06 nrd=1.14685 nrs=1.98347 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=26050 $Y=27490 $D=28
M4665 4324 78 VSS VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.41292e-13 pd=9.2e-07 ps=1.37846e-06 nrd=0.321429 nrs=0.450549 sa=5.4e-07 sb=1.96e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=26570 $Y=27150 $D=28
M4666 83 4322 4324 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.008e-13 pd=9.2e-07 ps=9.2e-07 nrd=0.321429 nrs=0.321429 sa=1.02e-06 sb=1.48e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=27050 $Y=27150 $D=28
M4667 4323 101 83 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.456e-13 as=1.008e-13 pd=1.08e-06 ps=9.2e-07 nrd=0.464286 nrs=0.321429 sa=1.5e-06 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=27530 $Y=27150 $D=28
M4668 VSS 4324 4323 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.52e-13 as=1.456e-13 pd=2.06667e-06 ps=1.08e-06 nrd=0.803571 nrs=0.464286 sa=1.95143e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=28170 $Y=27150 $D=28
M4669 VSS 163 4325 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55077e-14 as=9.6e-14 pd=5.41538e-07 ps=1.28e-06 nrd=1.14685 nrs=1.98347 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=46850 $Y=32290 $D=28
M4670 4327 176 VSS VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.41292e-13 pd=9.2e-07 ps=1.37846e-06 nrd=0.321429 nrs=0.450549 sa=5.4e-07 sb=1.96e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=47370 $Y=32290 $D=28
M4671 164 4325 4327 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.008e-13 pd=9.2e-07 ps=9.2e-07 nrd=0.321429 nrs=0.321429 sa=1.02e-06 sb=1.48e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=47850 $Y=32290 $D=28
M4672 4326 163 164 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.456e-13 as=1.008e-13 pd=1.08e-06 ps=9.2e-07 nrd=0.464286 nrs=0.321429 sa=1.5e-06 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=48330 $Y=32290 $D=28
M4673 VSS 4327 4326 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.52e-13 as=1.456e-13 pd=2.06667e-06 ps=1.08e-06 nrd=0.803571 nrs=0.464286 sa=1.95143e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=48970 $Y=32290 $D=28
M4674 VSS 114 4328 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55077e-14 as=9.6e-14 pd=5.41538e-07 ps=1.28e-06 nrd=1.14685 nrs=1.98347 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=48850 $Y=49090 $D=28
M4675 4330 183 VSS VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.41292e-13 pd=9.2e-07 ps=1.37846e-06 nrd=0.321429 nrs=0.450549 sa=5.4e-07 sb=1.96e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=49370 $Y=48750 $D=28
M4676 185 4328 4330 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.008e-13 pd=9.2e-07 ps=9.2e-07 nrd=0.321429 nrs=0.321429 sa=1.02e-06 sb=1.48e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=49850 $Y=48750 $D=28
M4677 4329 114 185 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.456e-13 as=1.008e-13 pd=1.08e-06 ps=9.2e-07 nrd=0.464286 nrs=0.321429 sa=1.5e-06 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=50330 $Y=48750 $D=28
M4678 VSS 4330 4329 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.52e-13 as=1.456e-13 pd=2.06667e-06 ps=1.08e-06 nrd=0.803571 nrs=0.464286 sa=1.95143e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=50970 $Y=48750 $D=28
M4679 VSS 114 4331 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55077e-14 as=9.6e-14 pd=5.41538e-07 ps=1.28e-06 nrd=1.14685 nrs=1.98347 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=50050 $Y=56290 $D=28
M4680 4333 186 VSS VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.41292e-13 pd=9.2e-07 ps=1.37846e-06 nrd=0.321429 nrs=0.450549 sa=5.4e-07 sb=1.96e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=50570 $Y=55950 $D=28
M4681 200 4331 4333 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.008e-13 pd=9.2e-07 ps=9.2e-07 nrd=0.321429 nrs=0.321429 sa=1.02e-06 sb=1.48e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=51050 $Y=55950 $D=28
M4682 4332 114 200 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.456e-13 as=1.008e-13 pd=1.08e-06 ps=9.2e-07 nrd=0.464286 nrs=0.321429 sa=1.5e-06 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=51530 $Y=55950 $D=28
M4683 VSS 4333 4332 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.52e-13 as=1.456e-13 pd=2.06667e-06 ps=1.08e-06 nrd=0.803571 nrs=0.464286 sa=1.95143e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=52170 $Y=55950 $D=28
M4684 VSS 816 4334 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55077e-14 as=9.6e-14 pd=5.41538e-07 ps=1.28e-06 nrd=1.14685 nrs=1.98347 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=58050 $Y=20290 $D=28
M4685 4336 235 VSS VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.41292e-13 pd=9.2e-07 ps=1.37846e-06 nrd=0.321429 nrs=0.450549 sa=5.4e-07 sb=1.96e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=58570 $Y=19950 $D=28
M4686 817 4334 4336 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.008e-13 pd=9.2e-07 ps=9.2e-07 nrd=0.321429 nrs=0.321429 sa=1.02e-06 sb=1.48e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=59050 $Y=19950 $D=28
M4687 4335 816 817 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.456e-13 as=1.008e-13 pd=1.08e-06 ps=9.2e-07 nrd=0.464286 nrs=0.321429 sa=1.5e-06 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=59530 $Y=19950 $D=28
M4688 VSS 4336 4335 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.52e-13 as=1.456e-13 pd=2.06667e-06 ps=1.08e-06 nrd=0.803571 nrs=0.464286 sa=1.95143e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=60170 $Y=19950 $D=28
M4689 VSS 228 4337 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55077e-14 as=9.6e-14 pd=5.41538e-07 ps=1.28e-06 nrd=1.14685 nrs=1.98347 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=68050 $Y=49090 $D=28
M4690 4339 283 VSS VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.41292e-13 pd=9.2e-07 ps=1.37846e-06 nrd=0.321429 nrs=0.450549 sa=5.4e-07 sb=1.96e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=68570 $Y=48750 $D=28
M4691 255 4337 4339 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.008e-13 pd=9.2e-07 ps=9.2e-07 nrd=0.321429 nrs=0.321429 sa=1.02e-06 sb=1.48e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=69050 $Y=48750 $D=28
M4692 4338 228 255 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.456e-13 as=1.008e-13 pd=1.08e-06 ps=9.2e-07 nrd=0.464286 nrs=0.321429 sa=1.5e-06 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=69530 $Y=48750 $D=28
M4693 VSS 4339 4338 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.52e-13 as=1.456e-13 pd=2.06667e-06 ps=1.08e-06 nrd=0.803571 nrs=0.464286 sa=1.95143e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=70170 $Y=48750 $D=28
M4694 VSS 411 4340 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55077e-14 as=9.6e-14 pd=5.41538e-07 ps=1.28e-06 nrd=1.14685 nrs=1.98347 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=100050 $Y=63490 $D=28
M4695 4342 372 VSS VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.41292e-13 pd=9.2e-07 ps=1.37846e-06 nrd=0.321429 nrs=0.450549 sa=5.4e-07 sb=1.96e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=100570 $Y=63150 $D=28
M4696 370 4340 4342 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.008e-13 pd=9.2e-07 ps=9.2e-07 nrd=0.321429 nrs=0.321429 sa=1.02e-06 sb=1.48e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=101050 $Y=63150 $D=28
M4697 4341 411 370 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.456e-13 as=1.008e-13 pd=1.08e-06 ps=9.2e-07 nrd=0.464286 nrs=0.321429 sa=1.5e-06 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=101530 $Y=63150 $D=28
M4698 VSS 4342 4341 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.52e-13 as=1.456e-13 pd=2.06667e-06 ps=1.08e-06 nrd=0.803571 nrs=0.464286 sa=1.95143e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=102170 $Y=63150 $D=28
M4699 4343 73 VSS VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.206e-13 as=2.144e-13 pd=1.03e-06 ps=1.98e-06 nrd=0.268657 nrs=0.477612 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=23210 $Y=55840 $D=28
M4700 VSS 73 4343 VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46642e-13 as=1.206e-13 pd=1.11245e-06 ps=1.03e-06 nrd=0.326669 nrs=0.268657 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=23690 $Y=55840 $D=28
M4701 82 4343 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.01358e-13 pd=1.28e-06 ps=1.52755e-06 nrd=0.195652 nrs=0.2379 sa=1.04826e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=24210 $Y=55590 $D=28
M4702 VSS 4343 82 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.52826e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=24690 $Y=55590 $D=28
M4703 82 4343 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.80435e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=25170 $Y=55590 $D=28
M4704 VSS 4343 82 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=1.93478e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=25650 $Y=55590 $D=28
M4705 4344 98 VSS VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.206e-13 as=2.144e-13 pd=1.03e-06 ps=1.98e-06 nrd=0.268657 nrs=0.477612 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=23610 $Y=41440 $D=28
M4706 VSS 98 4344 VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46642e-13 as=1.206e-13 pd=1.11245e-06 ps=1.03e-06 nrd=0.326669 nrs=0.268657 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=24090 $Y=41440 $D=28
M4707 84 4344 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.01358e-13 pd=1.28e-06 ps=1.52755e-06 nrd=0.195652 nrs=0.2379 sa=1.04826e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=24610 $Y=41190 $D=28
M4708 VSS 4344 84 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.52826e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=25090 $Y=41190 $D=28
M4709 84 4344 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.80435e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=25570 $Y=41190 $D=28
M4710 VSS 4344 84 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=1.93478e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=26050 $Y=41190 $D=28
M4711 4345 114 VSS VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.206e-13 as=2.144e-13 pd=1.03e-06 ps=1.98e-06 nrd=0.268657 nrs=0.477612 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=31610 $Y=27040 $D=28
M4712 VSS 114 4345 VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46642e-13 as=1.206e-13 pd=1.11245e-06 ps=1.03e-06 nrd=0.326669 nrs=0.268657 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=32090 $Y=27040 $D=28
M4713 113 4345 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.01358e-13 pd=1.28e-06 ps=1.52755e-06 nrd=0.195652 nrs=0.2379 sa=1.04826e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=32610 $Y=26790 $D=28
M4714 VSS 4345 113 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.52826e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=33090 $Y=26790 $D=28
M4715 113 4345 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.80435e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=33570 $Y=26790 $D=28
M4716 VSS 4345 113 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=1.93478e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=34050 $Y=26790 $D=28
M4717 4346 111 VSS VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.206e-13 as=2.144e-13 pd=1.03e-06 ps=1.98e-06 nrd=0.268657 nrs=0.477612 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=33210 $Y=75490 $D=28
M4718 VSS 111 4346 VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46642e-13 as=1.206e-13 pd=1.11245e-06 ps=1.03e-06 nrd=0.326669 nrs=0.268657 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=33690 $Y=75490 $D=28
M4719 89 4346 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.01358e-13 pd=1.28e-06 ps=1.52755e-06 nrd=0.195652 nrs=0.2379 sa=1.04826e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=34210 $Y=75490 $D=28
M4720 VSS 4346 89 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.52826e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=34690 $Y=75490 $D=28
M4721 89 4346 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.80435e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=35170 $Y=75490 $D=28
M4722 VSS 4346 89 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=1.93478e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=35650 $Y=75490 $D=28
M4723 4347 136 VSS VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.206e-13 as=2.144e-13 pd=1.03e-06 ps=1.98e-06 nrd=0.268657 nrs=0.477612 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=37210 $Y=46690 $D=28
M4724 VSS 136 4347 VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46642e-13 as=1.206e-13 pd=1.11245e-06 ps=1.03e-06 nrd=0.326669 nrs=0.268657 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=37690 $Y=46690 $D=28
M4725 176 4347 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.01358e-13 pd=1.28e-06 ps=1.52755e-06 nrd=0.195652 nrs=0.2379 sa=1.04826e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=38210 $Y=46690 $D=28
M4726 VSS 4347 176 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.52826e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=38690 $Y=46690 $D=28
M4727 176 4347 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.80435e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=39170 $Y=46690 $D=28
M4728 VSS 4347 176 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=1.93478e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=39650 $Y=46690 $D=28
M4729 4348 129 VSS VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.206e-13 as=2.144e-13 pd=1.03e-06 ps=1.98e-06 nrd=0.268657 nrs=0.477612 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=49610 $Y=41440 $D=28
M4730 VSS 129 4348 VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46642e-13 as=1.206e-13 pd=1.11245e-06 ps=1.03e-06 nrd=0.326669 nrs=0.268657 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=50090 $Y=41440 $D=28
M4731 228 4348 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.01358e-13 pd=1.28e-06 ps=1.52755e-06 nrd=0.195652 nrs=0.2379 sa=1.04826e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=50610 $Y=41190 $D=28
M4732 VSS 4348 228 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.52826e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=51090 $Y=41190 $D=28
M4733 228 4348 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.80435e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=51570 $Y=41190 $D=28
M4734 VSS 4348 228 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=1.93478e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=52050 $Y=41190 $D=28
M4735 4349 283 VSS VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.206e-13 as=2.144e-13 pd=1.03e-06 ps=1.98e-06 nrd=0.268657 nrs=0.477612 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=75610 $Y=46690 $D=28
M4736 VSS 283 4349 VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46642e-13 as=1.206e-13 pd=1.11245e-06 ps=1.03e-06 nrd=0.326669 nrs=0.268657 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=76090 $Y=46690 $D=28
M4737 354 4349 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.01358e-13 pd=1.28e-06 ps=1.52755e-06 nrd=0.195652 nrs=0.2379 sa=1.04826e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=76610 $Y=46690 $D=28
M4738 VSS 4349 354 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.52826e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=77090 $Y=46690 $D=28
M4739 354 4349 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.80435e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=77570 $Y=46690 $D=28
M4740 VSS 4349 354 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=1.93478e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=78050 $Y=46690 $D=28
M4741 4350 354 VSS VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.206e-13 as=2.144e-13 pd=1.03e-06 ps=1.98e-06 nrd=0.268657 nrs=0.477612 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=98810 $Y=48640 $D=28
M4742 VSS 354 4350 VSS lpnfet w=6.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46642e-13 as=1.206e-13 pd=1.11245e-06 ps=1.03e-06 nrd=0.326669 nrs=0.268657 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.04e-14 panw9=0 panw10=0 $X=99290 $Y=48640 $D=28
M4743 395 4350 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.01358e-13 pd=1.28e-06 ps=1.52755e-06 nrd=0.195652 nrs=0.2379 sa=1.04826e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=99810 $Y=48390 $D=28
M4744 VSS 4350 395 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.52826e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=100290 $Y=48390 $D=28
M4745 395 4350 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=1.656e-13 pd=1.28e-06 ps=1.28e-06 nrd=0.195652 nrs=0.195652 sa=1.80435e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=100770 $Y=48390 $D=28
M4746 VSS 4350 395 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=1.93478e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=101250 $Y=48390 $D=28
M4747 4351 86 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=28630 $Y=55960 $D=28
M4748 VSS 86 4351 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26612e-13 as=9.9e-14 pd=9.87755e-07 ps=9.1e-07 nrd=0.418553 nrs=0.327273 sa=8e-07 sb=1.88e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=29110 $Y=55960 $D=28
M4749 114 4351 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.11788e-13 pd=1.28e-06 ps=1.65224e-06 nrd=0.195652 nrs=0.250222 sa=9.17826e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=29630 $Y=55590 $D=28
M4750 VSS 4351 114 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=1.39783e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=30110 $Y=55590 $D=28
M4751 114 4351 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.08475e-13 pd=2.48e-06 ps=1.41472e-06 nrd=0.347826 nrs=0.246308 sa=1.74261e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=30670 $Y=55590 $D=28
M4752 4352 89 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=30230 $Y=75490 $D=28
M4753 VSS 89 4352 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26612e-13 as=9.9e-14 pd=9.87755e-07 ps=9.1e-07 nrd=0.418553 nrs=0.327273 sa=8e-07 sb=1.88e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=30710 $Y=75490 $D=28
M4754 162 4352 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.11788e-13 pd=1.28e-06 ps=1.65224e-06 nrd=0.195652 nrs=0.250222 sa=9.17826e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=31230 $Y=75490 $D=28
M4755 VSS 4352 162 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=1.39783e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=31710 $Y=75490 $D=28
M4756 162 4352 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.08475e-13 pd=2.48e-06 ps=1.41472e-06 nrd=0.347826 nrs=0.246308 sa=1.74261e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=32270 $Y=75490 $D=28
M4757 4353 114 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=37030 $Y=48760 $D=28
M4758 VSS 114 4353 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26612e-13 as=9.9e-14 pd=9.87755e-07 ps=9.1e-07 nrd=0.418553 nrs=0.327273 sa=8e-07 sb=1.88e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=37510 $Y=48760 $D=28
M4759 163 4353 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.11788e-13 pd=1.28e-06 ps=1.65224e-06 nrd=0.195652 nrs=0.250222 sa=9.17826e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=38030 $Y=48390 $D=28
M4760 VSS 4353 163 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=1.39783e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=38510 $Y=48390 $D=28
M4761 163 4353 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.08475e-13 pd=2.48e-06 ps=1.41472e-06 nrd=0.347826 nrs=0.246308 sa=1.74261e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=39070 $Y=48390 $D=28
M4762 4354 894 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=48230 $Y=63160 $D=28
M4763 VSS 894 4354 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26612e-13 as=9.9e-14 pd=9.87755e-07 ps=9.1e-07 nrd=0.418553 nrs=0.327273 sa=8e-07 sb=1.88e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=48710 $Y=63160 $D=28
M4764 248 4354 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.11788e-13 pd=1.28e-06 ps=1.65224e-06 nrd=0.195652 nrs=0.250222 sa=9.17826e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=49230 $Y=62790 $D=28
M4765 VSS 4354 248 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=1.39783e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=49710 $Y=62790 $D=28
M4766 248 4354 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.08475e-13 pd=2.48e-06 ps=1.41472e-06 nrd=0.347826 nrs=0.246308 sa=1.74261e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=50270 $Y=62790 $D=28
M4767 4355 182 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=49430 $Y=25090 $D=28
M4768 VSS 182 4355 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26612e-13 as=9.9e-14 pd=9.87755e-07 ps=9.1e-07 nrd=0.418553 nrs=0.327273 sa=8e-07 sb=1.88e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=49910 $Y=25090 $D=28
M4769 198 4355 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.11788e-13 pd=1.28e-06 ps=1.65224e-06 nrd=0.195652 nrs=0.250222 sa=9.17826e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=50430 $Y=25090 $D=28
M4770 VSS 4355 198 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=1.39783e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=50910 $Y=25090 $D=28
M4771 198 4355 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.08475e-13 pd=2.48e-06 ps=1.41472e-06 nrd=0.347826 nrs=0.246308 sa=1.74261e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=51470 $Y=25090 $D=28
M4772 4356 213 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=71430 $Y=48760 $D=28
M4773 VSS 213 4356 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26612e-13 as=9.9e-14 pd=9.87755e-07 ps=9.1e-07 nrd=0.418553 nrs=0.327273 sa=8e-07 sb=1.88e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=71910 $Y=48760 $D=28
M4774 325 4356 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.11788e-13 pd=1.28e-06 ps=1.65224e-06 nrd=0.195652 nrs=0.250222 sa=9.17826e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=72430 $Y=48390 $D=28
M4775 VSS 4356 325 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=1.39783e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=72910 $Y=48390 $D=28
M4776 325 4356 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.08475e-13 pd=2.48e-06 ps=1.41472e-06 nrd=0.347826 nrs=0.246308 sa=1.74261e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=73470 $Y=48390 $D=28
M4777 4357 320 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=81030 $Y=48760 $D=28
M4778 VSS 320 4357 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26612e-13 as=9.9e-14 pd=9.87755e-07 ps=9.1e-07 nrd=0.418553 nrs=0.327273 sa=8e-07 sb=1.88e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=81510 $Y=48760 $D=28
M4779 311 4357 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.11788e-13 pd=1.28e-06 ps=1.65224e-06 nrd=0.195652 nrs=0.250222 sa=9.17826e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=82030 $Y=48390 $D=28
M4780 VSS 4357 311 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=1.39783e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=82510 $Y=48390 $D=28
M4781 311 4357 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.08475e-13 pd=2.48e-06 ps=1.41472e-06 nrd=0.347826 nrs=0.246308 sa=1.74261e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=83070 $Y=48390 $D=28
M4782 4358 346 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=83030 $Y=39490 $D=28
M4783 VSS 346 4358 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26612e-13 as=9.9e-14 pd=9.87755e-07 ps=9.1e-07 nrd=0.418553 nrs=0.327273 sa=8e-07 sb=1.88e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=83510 $Y=39490 $D=28
M4784 350 4358 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.11788e-13 pd=1.28e-06 ps=1.65224e-06 nrd=0.195652 nrs=0.250222 sa=9.17826e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=84030 $Y=39490 $D=28
M4785 VSS 4358 350 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=1.39783e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=84510 $Y=39490 $D=28
M4786 350 4358 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.08475e-13 pd=2.48e-06 ps=1.41472e-06 nrd=0.347826 nrs=0.246308 sa=1.74261e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=85070 $Y=39490 $D=28
M4787 4359 325 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=89830 $Y=46690 $D=28
M4788 VSS 325 4359 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26612e-13 as=9.9e-14 pd=9.87755e-07 ps=9.1e-07 nrd=0.418553 nrs=0.327273 sa=8e-07 sb=1.88e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=90310 $Y=46690 $D=28
M4789 400 4359 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.11788e-13 pd=1.28e-06 ps=1.65224e-06 nrd=0.195652 nrs=0.250222 sa=9.17826e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=90830 $Y=46690 $D=28
M4790 VSS 4359 400 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=1.39783e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=91310 $Y=46690 $D=28
M4791 400 4359 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.08475e-13 pd=2.48e-06 ps=1.41472e-06 nrd=0.347826 nrs=0.246308 sa=1.74261e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=91870 $Y=46690 $D=28
M4792 4360 246 VSS VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.9e-14 as=1.76e-13 pd=9.1e-07 ps=1.74e-06 nrd=0.327273 nrs=0.581818 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=93030 $Y=46690 $D=28
M4793 VSS 246 4360 VSS lpnfet w=5.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26612e-13 as=9.9e-14 pd=9.87755e-07 ps=9.1e-07 nrd=0.418553 nrs=0.327273 sa=8e-07 sb=1.88e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=93510 $Y=46690 $D=28
M4794 410 4360 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.11788e-13 pd=1.28e-06 ps=1.65224e-06 nrd=0.195652 nrs=0.250222 sa=9.17826e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=94030 $Y=46690 $D=28
M4795 VSS 4360 410 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.08475e-13 as=1.656e-13 pd=1.41472e-06 ps=1.28e-06 nrd=0.246308 nrs=0.195652 sa=1.39783e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=94510 $Y=46690 $D=28
M4796 410 4360 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.08475e-13 pd=2.48e-06 ps=1.41472e-06 nrd=0.347826 nrs=0.246308 sa=1.74261e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=95070 $Y=46690 $D=28
M4797 291 284 VSS VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.36e-14 as=1.664e-13 pd=8.8e-07 ps=1.68e-06 nrd=0.346154 nrs=0.615385 sa=3.2e-07 sb=1.22e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=76010 $Y=34390 $D=28
M4798 VSS 284 291 VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.78563e-13 as=9.36e-14 pd=1.43661e-06 ps=8.8e-07 nrd=0.660365 nrs=0.346154 sa=8e-07 sb=7.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=76490 $Y=34390 $D=28
M4799 291 284 VSS VSS lpnfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.216e-13 as=1.30488e-13 pd=1.4e-06 ps=1.04983e-06 nrd=0.842105 nrs=0.903657 sa=1.36e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=9.6e-15 panw8=0 panw9=0 panw10=0 $X=77050 $Y=34530 $D=28
M4800 304 284 VSS VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.36e-14 as=1.664e-13 pd=8.8e-07 ps=1.68e-06 nrd=0.346154 nrs=0.615385 sa=3.2e-07 sb=1.22e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=78010 $Y=34390 $D=28
M4801 VSS 284 304 VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.78563e-13 as=9.36e-14 pd=1.43661e-06 ps=8.8e-07 nrd=0.660365 nrs=0.346154 sa=8e-07 sb=7.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=78490 $Y=34390 $D=28
M4802 304 284 VSS VSS lpnfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.216e-13 as=1.30488e-13 pd=1.4e-06 ps=1.04983e-06 nrd=0.842105 nrs=0.903657 sa=1.36e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=9.6e-15 panw8=0 panw9=0 panw10=0 $X=79050 $Y=34530 $D=28
M4803 316 302 VSS VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.36e-14 as=1.664e-13 pd=8.8e-07 ps=1.68e-06 nrd=0.346154 nrs=0.615385 sa=3.2e-07 sb=1.22e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=84010 $Y=12790 $D=28
M4804 VSS 302 316 VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.78563e-13 as=9.36e-14 pd=1.43661e-06 ps=8.8e-07 nrd=0.660365 nrs=0.346154 sa=8e-07 sb=7.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=84490 $Y=12790 $D=28
M4805 316 302 VSS VSS lpnfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.216e-13 as=1.30488e-13 pd=1.4e-06 ps=1.04983e-06 nrd=0.842105 nrs=0.903657 sa=1.36e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=9.6e-15 panw8=0 panw9=0 panw10=0 $X=85050 $Y=12930 $D=28
M4806 265 242 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.004e-13 as=1.004e-13 pd=1.3e-06 ps=1.3e-06 nrd=1.74306 nrs=1.74306 sa=3.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=68570 $Y=46690 $D=28
M4807 297 313 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.004e-13 as=1.004e-13 pd=1.3e-06 ps=1.3e-06 nrd=1.74306 nrs=1.74306 sa=3.6e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=4.8e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=78570 $Y=41870 $D=28
M4808 4369 4361 4362 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=12860 $Y=13090 $D=28
M4809 4371 798 4369 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=13180 $Y=13090 $D=28
M4810 VSS 76 4371 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=13500 $Y=13090 $D=28
M4811 VSS clk 4361 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=14480 $Y=12840 $D=28
M4812 4364 4361 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.084e-13 as=7.56667e-14 pd=1.38e-06 ps=7.48718e-07 nrd=2.71 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=14990 $Y=12940 $D=28
M4813 4373 4364 4362 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.608e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=16010 $Y=13010 $D=28
M4814 4374 4363 4373 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=1.288e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=16330 $Y=13010 $D=28
M4815 VSS 76 4374 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.052e-13 as=2e-14 pd=1.3e-06 ps=4e-07 nrd=2.63 nrs=0.5 sa=1e-06 sb=9.68e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=16650 $Y=13010 $D=28
M4816 4363 4362 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.88e-14 as=1.052e-13 pd=9.6e-07 ps=1.3e-06 nrd=2.22 nrs=2.63 sa=1.44e-06 sb=5.28e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=17090 $Y=13010 $D=28
M4817 4365 4364 4363 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76e-14 as=8.88e-14 pd=8.8e-07 ps=9.6e-07 nrd=1.94 nrs=2.22 sa=8.52e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=3.6e-15 panw8=2.04e-14 panw9=0 panw10=0 $X=17650 $Y=12870 $D=28
M4818 4376 4361 4365 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=7.76e-14 pd=4e-07 ps=8.8e-07 nrd=0.5 nrs=1.94 sa=3.6e-07 sb=1.42e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=18210 $Y=13110 $D=28
M4819 VSS 4368 4376 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13103e-14 as=2e-14 pd=4.72414e-07 ps=4e-07 nrd=1.53276 nrs=0.5 sa=6.8e-07 sb=1.1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=18530 $Y=13110 $D=28
M4820 4377 76 VSS VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.2e-14 as=1.59407e-13 pd=7.2e-07 ps=1.22828e-06 nrd=0.192308 nrs=0.589523 sa=5.83077e-07 sb=6.04615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=18970 $Y=12790 $D=28
M4821 4368 4365 4377 VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48e-13 as=5.2e-14 pd=1.72e-06 ps=7.2e-07 nrd=0.547337 nrs=0.192308 sa=9.03077e-07 sb=2.84615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=19290 $Y=12790 $D=28
M4822 4366 4368 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=6.74414e-14 pd=1.28e-06 ps=5.19655e-07 nrd=1.98347 nrs=1.39342 sa=5.58182e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.64e-14 panw10=0 $X=19730 $Y=12390 $D=28
M4823 VSS 4366 4367 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.368e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.279773 sa=2.57391e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=20590 $Y=12390 $D=28
M4824 62 4368 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=7.37391e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=21070 $Y=12390 $D=28
M4825 4386 4378 4379 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=16060 $Y=61110 $D=28
M4826 4388 24 4386 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=16380 $Y=61110 $D=28
M4827 VSS 32 4388 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=16700 $Y=61110 $D=28
M4828 VSS clk 4378 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=17680 $Y=61260 $D=28
M4829 4381 4378 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.084e-13 as=7.56667e-14 pd=1.38e-06 ps=7.48718e-07 nrd=2.71 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=18190 $Y=61260 $D=28
M4830 4390 4381 4379 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.608e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=19210 $Y=61190 $D=28
M4831 4391 4380 4390 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=1.288e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=19530 $Y=61190 $D=28
M4832 VSS 32 4391 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.052e-13 as=2e-14 pd=1.3e-06 ps=4e-07 nrd=2.63 nrs=0.5 sa=1e-06 sb=9.68e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=19850 $Y=61190 $D=28
M4833 4380 4379 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.88e-14 as=1.052e-13 pd=9.6e-07 ps=1.3e-06 nrd=2.22 nrs=2.63 sa=1.44e-06 sb=5.28e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=20290 $Y=61190 $D=28
M4834 4382 4381 4380 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76e-14 as=8.88e-14 pd=8.8e-07 ps=9.6e-07 nrd=1.94 nrs=2.22 sa=8.52e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=3.6e-15 panw8=2.04e-14 panw9=0 panw10=0 $X=20850 $Y=61330 $D=28
M4835 4393 4378 4382 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=7.76e-14 pd=4e-07 ps=8.8e-07 nrd=0.5 nrs=1.94 sa=3.6e-07 sb=1.42e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=21410 $Y=61090 $D=28
M4836 VSS 4385 4393 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13103e-14 as=2e-14 pd=4.72414e-07 ps=4e-07 nrd=1.53276 nrs=0.5 sa=6.8e-07 sb=1.1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=21730 $Y=61090 $D=28
M4837 4394 32 VSS VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.2e-14 as=1.59407e-13 pd=7.2e-07 ps=1.22828e-06 nrd=0.192308 nrs=0.589523 sa=5.83077e-07 sb=6.04615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=22170 $Y=61090 $D=28
M4838 4385 4382 4394 VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48e-13 as=5.2e-14 pd=1.72e-06 ps=7.2e-07 nrd=0.547337 nrs=0.192308 sa=9.03077e-07 sb=2.84615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=22490 $Y=61090 $D=28
M4839 4383 4385 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=6.74414e-14 pd=1.28e-06 ps=5.19655e-07 nrd=1.98347 nrs=1.39342 sa=5.58182e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.64e-14 panw10=0 $X=22930 $Y=61790 $D=28
M4840 VSS 4383 4384 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.368e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.279773 sa=2.57391e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=23790 $Y=61090 $D=28
M4841 109 4385 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=7.37391e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=24270 $Y=61090 $D=28
M4842 4403 4395 4396 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=16860 $Y=39510 $D=28
M4843 4405 801 4403 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=17180 $Y=39510 $D=28
M4844 VSS 68 4405 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=17500 $Y=39510 $D=28
M4845 VSS clk 4395 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=18480 $Y=39660 $D=28
M4846 4398 4395 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.084e-13 as=7.56667e-14 pd=1.38e-06 ps=7.48718e-07 nrd=2.71 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=18990 $Y=39660 $D=28
M4847 4407 4398 4396 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.608e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=20010 $Y=39590 $D=28
M4848 4408 4397 4407 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=1.288e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=20330 $Y=39590 $D=28
M4849 VSS 68 4408 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.052e-13 as=2e-14 pd=1.3e-06 ps=4e-07 nrd=2.63 nrs=0.5 sa=1e-06 sb=9.68e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=20650 $Y=39590 $D=28
M4850 4397 4396 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.88e-14 as=1.052e-13 pd=9.6e-07 ps=1.3e-06 nrd=2.22 nrs=2.63 sa=1.44e-06 sb=5.28e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=21090 $Y=39590 $D=28
M4851 4399 4398 4397 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76e-14 as=8.88e-14 pd=8.8e-07 ps=9.6e-07 nrd=1.94 nrs=2.22 sa=8.52e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=3.6e-15 panw8=2.04e-14 panw9=0 panw10=0 $X=21650 $Y=39730 $D=28
M4852 4410 4395 4399 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=7.76e-14 pd=4e-07 ps=8.8e-07 nrd=0.5 nrs=1.94 sa=3.6e-07 sb=1.42e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=22210 $Y=39490 $D=28
M4853 VSS 4402 4410 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13103e-14 as=2e-14 pd=4.72414e-07 ps=4e-07 nrd=1.53276 nrs=0.5 sa=6.8e-07 sb=1.1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=22530 $Y=39490 $D=28
M4854 4411 68 VSS VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.2e-14 as=1.59407e-13 pd=7.2e-07 ps=1.22828e-06 nrd=0.192308 nrs=0.589523 sa=5.83077e-07 sb=6.04615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=22970 $Y=39490 $D=28
M4855 4402 4399 4411 VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48e-13 as=5.2e-14 pd=1.72e-06 ps=7.2e-07 nrd=0.547337 nrs=0.192308 sa=9.03077e-07 sb=2.84615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=23290 $Y=39490 $D=28
M4856 4400 4402 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=6.74414e-14 pd=1.28e-06 ps=5.19655e-07 nrd=1.98347 nrs=1.39342 sa=5.58182e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.64e-14 panw10=0 $X=23730 $Y=40190 $D=28
M4857 VSS 4400 4401 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.368e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.279773 sa=2.57391e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=24590 $Y=39490 $D=28
M4858 159 4402 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=7.37391e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=25070 $Y=39490 $D=28
M4859 4420 4412 4413 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=54460 $Y=13090 $D=28
M4860 4422 226 4420 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=54780 $Y=13090 $D=28
M4861 VSS 202 4422 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=55100 $Y=13090 $D=28
M4862 VSS clk 4412 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=56080 $Y=12840 $D=28
M4863 4415 4412 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.084e-13 as=7.56667e-14 pd=1.38e-06 ps=7.48718e-07 nrd=2.71 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=56590 $Y=12940 $D=28
M4864 4424 4415 4413 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.608e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=57610 $Y=13010 $D=28
M4865 4425 4414 4424 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=1.288e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=57930 $Y=13010 $D=28
M4866 VSS 202 4425 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.052e-13 as=2e-14 pd=1.3e-06 ps=4e-07 nrd=2.63 nrs=0.5 sa=1e-06 sb=9.68e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=58250 $Y=13010 $D=28
M4867 4414 4413 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.88e-14 as=1.052e-13 pd=9.6e-07 ps=1.3e-06 nrd=2.22 nrs=2.63 sa=1.44e-06 sb=5.28e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=58690 $Y=13010 $D=28
M4868 4416 4415 4414 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76e-14 as=8.88e-14 pd=8.8e-07 ps=9.6e-07 nrd=1.94 nrs=2.22 sa=8.52e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=3.6e-15 panw8=2.04e-14 panw9=0 panw10=0 $X=59250 $Y=12870 $D=28
M4869 4427 4412 4416 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=7.76e-14 pd=4e-07 ps=8.8e-07 nrd=0.5 nrs=1.94 sa=3.6e-07 sb=1.42e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=59810 $Y=13110 $D=28
M4870 VSS 4419 4427 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13103e-14 as=2e-14 pd=4.72414e-07 ps=4e-07 nrd=1.53276 nrs=0.5 sa=6.8e-07 sb=1.1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=60130 $Y=13110 $D=28
M4871 4428 202 VSS VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.2e-14 as=1.59407e-13 pd=7.2e-07 ps=1.22828e-06 nrd=0.192308 nrs=0.589523 sa=5.83077e-07 sb=6.04615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=60570 $Y=12790 $D=28
M4872 4419 4416 4428 VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48e-13 as=5.2e-14 pd=1.72e-06 ps=7.2e-07 nrd=0.547337 nrs=0.192308 sa=9.03077e-07 sb=2.84615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=60890 $Y=12790 $D=28
M4873 4417 4419 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=6.74414e-14 pd=1.28e-06 ps=5.19655e-07 nrd=1.98347 nrs=1.39342 sa=5.58182e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.64e-14 panw10=0 $X=61330 $Y=12390 $D=28
M4874 VSS 4417 4418 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.368e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.279773 sa=2.57391e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=62190 $Y=12390 $D=28
M4875 143 4419 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=7.37391e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=62670 $Y=12390 $D=28
M4876 4437 4429 4430 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=62860 $Y=17910 $D=28
M4877 4439 261 4437 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=63180 $Y=17910 $D=28
M4878 VSS 299 4439 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=63500 $Y=17910 $D=28
M4879 VSS clk 4429 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=64480 $Y=18060 $D=28
M4880 4432 4429 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.084e-13 as=7.56667e-14 pd=1.38e-06 ps=7.48718e-07 nrd=2.71 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=64990 $Y=18060 $D=28
M4881 4441 4432 4430 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.608e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=66010 $Y=17990 $D=28
M4882 4442 4431 4441 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=1.288e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=66330 $Y=17990 $D=28
M4883 VSS 299 4442 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.052e-13 as=2e-14 pd=1.3e-06 ps=4e-07 nrd=2.63 nrs=0.5 sa=1e-06 sb=9.68e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=66650 $Y=17990 $D=28
M4884 4431 4430 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.88e-14 as=1.052e-13 pd=9.6e-07 ps=1.3e-06 nrd=2.22 nrs=2.63 sa=1.44e-06 sb=5.28e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=67090 $Y=17990 $D=28
M4885 4433 4432 4431 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76e-14 as=8.88e-14 pd=8.8e-07 ps=9.6e-07 nrd=1.94 nrs=2.22 sa=8.52e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=3.6e-15 panw8=2.04e-14 panw9=0 panw10=0 $X=67650 $Y=18130 $D=28
M4886 4444 4429 4433 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=7.76e-14 pd=4e-07 ps=8.8e-07 nrd=0.5 nrs=1.94 sa=3.6e-07 sb=1.42e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=68210 $Y=17890 $D=28
M4887 VSS 4436 4444 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13103e-14 as=2e-14 pd=4.72414e-07 ps=4e-07 nrd=1.53276 nrs=0.5 sa=6.8e-07 sb=1.1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=68530 $Y=17890 $D=28
M4888 4445 299 VSS VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.2e-14 as=1.59407e-13 pd=7.2e-07 ps=1.22828e-06 nrd=0.192308 nrs=0.589523 sa=5.83077e-07 sb=6.04615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=68970 $Y=17890 $D=28
M4889 4436 4433 4445 VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48e-13 as=5.2e-14 pd=1.72e-06 ps=7.2e-07 nrd=0.547337 nrs=0.192308 sa=9.03077e-07 sb=2.84615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=69290 $Y=17890 $D=28
M4890 4434 4436 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=6.74414e-14 pd=1.28e-06 ps=5.19655e-07 nrd=1.98347 nrs=1.39342 sa=5.58182e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.64e-14 panw10=0 $X=69730 $Y=18590 $D=28
M4891 VSS 4434 4435 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.368e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.279773 sa=2.57391e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=70590 $Y=17890 $D=28
M4892 264 4436 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=7.37391e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=71070 $Y=17890 $D=28
M4893 4454 4446 4447 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=1.272e-13 pd=4e-07 ps=1.52e-06 nrd=0.5 nrs=3.18 sa=3.7e-07 sb=1e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=77260 $Y=25110 $D=28
M4894 4456 827 4454 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.9e-07 sb=6.8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=77580 $Y=25110 $D=28
M4895 VSS 303 4456 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.43167e-13 as=2e-14 pd=1.275e-06 ps=4e-07 nrd=3.57917 nrs=0.5 sa=1.01e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=2.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=77900 $Y=25110 $D=28
M4896 VSS clk 4446 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.135e-13 as=9.6e-14 pd=1.12308e-06 ps=1.24e-06 nrd=1.26111 nrs=1.06667 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=2.04e-14 panw8=0 panw9=0 panw10=0 $X=78880 $Y=25260 $D=28
M4897 4449 4446 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.084e-13 as=7.56667e-14 pd=1.38e-06 ps=7.48718e-07 nrd=2.71 nrs=1.89167 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.6e-15 panw6=1.2e-14 panw7=8.4e-15 panw8=0 panw9=0 panw10=0 $X=79390 $Y=25260 $D=28
M4898 4458 4449 4447 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=9.72e-14 pd=4e-07 ps=1.3e-06 nrd=0.5 nrs=2.43 sa=3.6e-07 sb=1.608e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=80410 $Y=25190 $D=28
M4899 4459 4448 4458 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=2e-14 pd=4e-07 ps=4e-07 nrd=0.5 nrs=0.5 sa=6.8e-07 sb=1.288e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=80730 $Y=25190 $D=28
M4900 VSS 303 4459 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.052e-13 as=2e-14 pd=1.3e-06 ps=4e-07 nrd=2.63 nrs=0.5 sa=1e-06 sb=9.68e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=81050 $Y=25190 $D=28
M4901 4448 4447 VSS VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.88e-14 as=1.052e-13 pd=9.6e-07 ps=1.3e-06 nrd=2.22 nrs=2.63 sa=1.44e-06 sb=5.28e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=81490 $Y=25190 $D=28
M4902 4450 4449 4448 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76e-14 as=8.88e-14 pd=8.8e-07 ps=9.6e-07 nrd=1.94 nrs=2.22 sa=8.52e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=3.6e-15 panw8=2.04e-14 panw9=0 panw10=0 $X=82050 $Y=25330 $D=28
M4903 4461 4446 4450 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2e-14 as=7.76e-14 pd=4e-07 ps=8.8e-07 nrd=0.5 nrs=1.94 sa=3.6e-07 sb=1.42e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=82610 $Y=25090 $D=28
M4904 VSS 4453 4461 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.13103e-14 as=2e-14 pd=4.72414e-07 ps=4e-07 nrd=1.53276 nrs=0.5 sa=6.8e-07 sb=1.1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 $X=82930 $Y=25090 $D=28
M4905 4462 303 VSS VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.2e-14 as=1.59407e-13 pd=7.2e-07 ps=1.22828e-06 nrd=0.192308 nrs=0.589523 sa=5.83077e-07 sb=6.04615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=83370 $Y=25090 $D=28
M4906 4453 4450 4462 VSS lpnfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.48e-13 as=5.2e-14 pd=1.72e-06 ps=7.2e-07 nrd=0.547337 nrs=0.192308 sa=9.03077e-07 sb=2.84615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=83690 $Y=25090 $D=28
M4907 4451 4453 VSS VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=6.74414e-14 pd=1.28e-06 ps=5.19655e-07 nrd=1.98347 nrs=1.39342 sa=5.58182e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=2.64e-14 panw10=0 $X=84130 $Y=25790 $D=28
M4908 VSS 4451 4452 VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.656e-13 as=2.368e-13 pd=1.28e-06 ps=2.48e-06 nrd=0.195652 nrs=0.279773 sa=2.57391e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=84990 $Y=25090 $D=28
M4909 298 4453 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.656e-13 pd=2.48e-06 ps=1.28e-06 nrd=0.347826 nrs=0.195652 sa=7.37391e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=85470 $Y=25090 $D=28
M4910 4464 22 4463 VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.604e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.369048 sa=3.1e-07 sb=1.825e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=12740 $Y=32290 $D=28
M4911 VSS 42 4464 VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.56361e-13 as=8.4e-14 pd=1.29542e-06 ps=1.04e-06 nrd=0.221601 nrs=0.119048 sa=6.3e-07 sb=1.7869e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=13060 $Y=32290 $D=28
M4912 4465 62 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.52639e-13 pd=1.02e-06 ps=1.26458e-06 nrd=0.121951 nrs=0.227006 sa=1.02683e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=13540 $Y=32390 $D=28
M4913 800 4463 4465 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.34683e-06 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=13860 $Y=32390 $D=28
M4914 4466 4463 800 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.82683e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=14340 $Y=32390 $D=28
M4915 VSS 62 4466 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.94049e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=14660 $Y=32390 $D=28
M4916 4467 62 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.98732e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=15140 $Y=32390 $D=28
M4917 800 4463 4467 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=15460 $Y=32390 $D=28
M4918 4469 215 4468 VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.604e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.369048 sa=3.1e-07 sb=1.825e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=59140 $Y=62870 $D=28
M4919 VSS 222 4469 VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.56361e-13 as=8.4e-14 pd=1.29542e-06 ps=1.04e-06 nrd=0.221601 nrs=0.119048 sa=6.3e-07 sb=1.7869e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=59460 $Y=62870 $D=28
M4920 4470 233 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.52639e-13 pd=1.02e-06 ps=1.26458e-06 nrd=0.121951 nrs=0.227006 sa=1.02683e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=59940 $Y=62790 $D=28
M4921 225 4468 4470 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.34683e-06 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=60260 $Y=62790 $D=28
M4922 4471 4468 225 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.82683e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=60740 $Y=62790 $D=28
M4923 VSS 233 4471 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.94049e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=61060 $Y=62790 $D=28
M4924 4472 233 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.98732e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=61540 $Y=62790 $D=28
M4925 225 4468 4472 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=61860 $Y=62790 $D=28
M4926 4474 265 4473 VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.604e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.369048 sa=3.1e-07 sb=1.825e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=71940 $Y=41270 $D=28
M4927 VSS 270 4474 VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.56361e-13 as=8.4e-14 pd=1.29542e-06 ps=1.04e-06 nrd=0.221601 nrs=0.119048 sa=6.3e-07 sb=1.7869e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=72260 $Y=41270 $D=28
M4928 4475 292 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.52639e-13 pd=1.02e-06 ps=1.26458e-06 nrd=0.121951 nrs=0.227006 sa=1.02683e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=72740 $Y=41190 $D=28
M4929 824 4473 4475 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.34683e-06 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=73060 $Y=41190 $D=28
M4930 4476 4473 824 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.82683e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=73540 $Y=41190 $D=28
M4931 VSS 292 4476 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.94049e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=73860 $Y=41190 $D=28
M4932 4477 292 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.98732e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=74340 $Y=41190 $D=28
M4933 824 4473 4477 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=8.2e-14 pd=2.28e-06 ps=1.02e-06 nrd=0.390244 nrs=0.121951 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=74660 $Y=41190 $D=28
M4934 VSS 45 4478 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.76632e-14 as=9.6e-14 pd=5.67368e-07 ps=1.28e-06 nrd=1.19139 nrs=1.98347 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=8.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=12850 $Y=56240 $D=28
M4935 4480 31 VSS VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.72e-14 as=1.41537e-13 pd=9e-07 ps=1.39263e-06 nrd=0.333333 nrs=0.48538 sa=5.64444e-07 sb=1.98e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=13410 $Y=55920 $D=28
M4936 25 45 4480 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.79855e-14 as=9.72e-14 pd=9.03273e-07 ps=9e-07 nrd=0.336027 nrs=0.333333 sa=1.04444e-06 sb=1.5e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=13890 $Y=55920 $D=28
M4937 4479 4478 25 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.01615e-13 pd=1.1e-06 ps=9.36727e-07 nrd=0.482143 nrs=0.324026 sa=1.47929e-06 sb=1.02e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=14370 $Y=55910 $D=28
M4938 VSS 4480 4479 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.44533e-13 as=1.512e-13 pd=2.01333e-06 ps=1.1e-06 nrd=0.779762 nrs=0.482143 sa=1.92714e-06 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=15030 $Y=55910 $D=28
M4939 VSS 192 4481 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.76632e-14 as=9.6e-14 pd=5.67368e-07 ps=1.28e-06 nrd=1.19139 nrs=1.98347 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=8.4e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=67250 $Y=34640 $D=28
M4940 4483 231 VSS VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.72e-14 as=1.41537e-13 pd=9e-07 ps=1.39263e-06 nrd=0.333333 nrs=0.48538 sa=5.64444e-07 sb=1.98e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=67810 $Y=34320 $D=28
M4941 820 192 4483 VSS lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.79855e-14 as=9.72e-14 pd=9.03273e-07 ps=9e-07 nrd=0.336027 nrs=0.333333 sa=1.04444e-06 sb=1.5e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.08e-14 panw9=0 panw10=0 $X=68290 $Y=34320 $D=28
M4942 4482 4481 820 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.01615e-13 pd=1.1e-06 ps=9.36727e-07 nrd=0.482143 nrs=0.324026 sa=1.47929e-06 sb=1.02e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=68770 $Y=34310 $D=28
M4943 VSS 4483 4482 VSS lpnfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.44533e-13 as=1.512e-13 pd=2.01333e-06 ps=1.1e-06 nrd=0.779762 nrs=0.482143 sa=1.92714e-06 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=69430 $Y=34310 $D=28
M4944 VSS 60 4484 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.15e-14 as=9.44e-14 pd=6.91667e-07 ps=1.28e-06 nrd=1.5375 nrs=2.36 sa=3.6e-07 sb=1.422e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=14960 $Y=68550 $D=28
M4945 4486 54 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.61e-14 pd=9.2e-07 ps=9.68333e-07 nrd=1.14286 nrs=1.09821 sa=7.6e-07 sb=7.47143e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=15520 $Y=68550 $D=28
M4946 41 60 4486 VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.59556e-14 as=8.96e-14 pd=7.67407e-07 ps=9.2e-07 nrd=0.84127 nrs=1.14286 sa=7.67143e-07 sb=9e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=16100 $Y=68370 $D=28
M4947 4485 4484 41 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.03037e-13 as=6.12444e-14 pd=1.01111e-06 ps=7.12593e-07 nrd=1.52422 nrs=0.905983 sa=1.26615e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=16680 $Y=68370 $D=28
M4948 VSS 4486 4485 VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.2e-14 as=1.10963e-13 pd=5.8e-07 ps=1.08889e-06 nrd=0.535714 nrs=1.41534 sa=6.9e-07 sb=7.22857e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=16880 $Y=69060 $D=28
M4949 VSS 116 4487 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.15e-14 as=9.44e-14 pd=6.91667e-07 ps=1.28e-06 nrd=1.5375 nrs=2.36 sa=3.6e-07 sb=1.422e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=34160 $Y=18150 $D=28
M4950 4489 118 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.61e-14 pd=9.2e-07 ps=9.68333e-07 nrd=1.14286 nrs=1.09821 sa=7.6e-07 sb=7.47143e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=34720 $Y=18150 $D=28
M4951 122 116 4489 VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.59556e-14 as=8.96e-14 pd=7.67407e-07 ps=9.2e-07 nrd=0.84127 nrs=1.14286 sa=7.67143e-07 sb=9e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=35300 $Y=17970 $D=28
M4952 4488 4487 122 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.03037e-13 as=6.12444e-14 pd=1.01111e-06 ps=7.12593e-07 nrd=1.52422 nrs=0.905983 sa=1.26615e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=35880 $Y=17970 $D=28
M4953 VSS 4489 4488 VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.2e-14 as=1.10963e-13 pd=5.8e-07 ps=1.08889e-06 nrd=0.535714 nrs=1.41534 sa=6.9e-07 sb=6.67143e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=36080 $Y=18660 $D=28
M4954 VSS 259 4490 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.15e-14 as=9.44e-14 pd=6.91667e-07 ps=1.28e-06 nrd=1.5375 nrs=2.36 sa=3.6e-07 sb=1.422e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=66560 $Y=20050 $D=28
M4955 4492 281 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=8.61e-14 pd=9.2e-07 ps=9.68333e-07 nrd=1.14286 nrs=1.09821 sa=7.6e-07 sb=7.47143e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=67120 $Y=19970 $D=28
M4956 257 259 4492 VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.59556e-14 as=8.96e-14 pd=7.67407e-07 ps=9.2e-07 nrd=0.84127 nrs=1.14286 sa=7.67143e-07 sb=9e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=67700 $Y=20150 $D=28
M4957 4491 4490 257 VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.03037e-13 as=6.12444e-14 pd=1.01111e-06 ps=7.12593e-07 nrd=1.52422 nrs=0.905983 sa=1.26615e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=68280 $Y=20170 $D=28
M4958 4491 4492 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10963e-13 as=4.2e-14 pd=1.08889e-06 ps=5.8e-07 nrd=1.41534 nrs=0.535714 sa=1.25821e-06 sb=6.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=68480 $Y=19620 $D=28
M4959 VSS 39 4493 VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.51504e-13 as=2.688e-13 pd=1.21446e-06 ps=2.32e-06 nrd=0.214716 nrs=0.380952 sa=3.2e-07 sb=1.95738e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=16260 $Y=17890 $D=28
M4960 4494 46 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.47896e-13 pd=1.02e-06 ps=1.18554e-06 nrd=0.121951 nrs=0.219953 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=16740 $Y=17890 $D=28
M4961 29 4493 4494 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.12e-06 sb=1.95634e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=17060 $Y=17890 $D=28
M4962 4495 4493 29 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.6e-06 sb=1.47634e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=17540 $Y=17890 $D=28
M4963 VSS 46 4495 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.92e-06 sb=1.15634e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=17860 $Y=17890 $D=28
M4964 4496 46 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=6.76341e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=18340 $Y=17890 $D=28
M4965 29 4493 4496 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.922e-13 as=8.2e-14 pd=2.38e-06 ps=1.02e-06 nrd=0.434563 nrs=0.121951 sa=2e-06 sb=3.56341e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=18660 $Y=17890 $D=28
M4966 VSS 162 4497 VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.51504e-13 as=2.688e-13 pd=1.21446e-06 ps=2.32e-06 nrd=0.214716 nrs=0.380952 sa=3.2e-07 sb=1.95738e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=53460 $Y=41270 $D=28
M4967 4498 135 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.47896e-13 pd=1.02e-06 ps=1.18554e-06 nrd=0.121951 nrs=0.219953 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=53940 $Y=41290 $D=28
M4968 206 4497 4498 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.12e-06 sb=1.95634e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=54260 $Y=41290 $D=28
M4969 4499 4497 206 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.6e-06 sb=1.47634e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=54740 $Y=41290 $D=28
M4970 VSS 135 4499 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.92e-06 sb=1.15634e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=55060 $Y=41290 $D=28
M4971 4500 135 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=6.76341e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=55540 $Y=41290 $D=28
M4972 206 4497 4500 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.922e-13 as=8.2e-14 pd=2.38e-06 ps=1.02e-06 nrd=0.434563 nrs=0.121951 sa=2e-06 sb=3.56341e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=55860 $Y=41290 $D=28
M4973 VSS 205 4501 VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.51504e-13 as=2.688e-13 pd=1.21446e-06 ps=2.32e-06 nrd=0.214716 nrs=0.380952 sa=3.2e-07 sb=1.95738e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=54660 $Y=25090 $D=28
M4974 4502 204 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.47896e-13 pd=1.02e-06 ps=1.18554e-06 nrd=0.121951 nrs=0.219953 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=55140 $Y=25090 $D=28
M4975 207 4501 4502 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.12e-06 sb=1.95634e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=55460 $Y=25090 $D=28
M4976 4503 4501 207 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.6e-06 sb=1.47634e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=55940 $Y=25090 $D=28
M4977 VSS 204 4503 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.92e-06 sb=1.15634e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=56260 $Y=25090 $D=28
M4978 4504 204 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=6.76341e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=56740 $Y=25090 $D=28
M4979 207 4501 4504 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.922e-13 as=8.2e-14 pd=2.38e-06 ps=1.02e-06 nrd=0.434563 nrs=0.121951 sa=2e-06 sb=3.56341e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=57060 $Y=25090 $D=28
M4980 VSS 135 4505 VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.51504e-13 as=2.688e-13 pd=1.21446e-06 ps=2.32e-06 nrd=0.214716 nrs=0.380952 sa=3.2e-07 sb=1.95738e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=61460 $Y=41270 $D=28
M4981 4506 162 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.47896e-13 pd=1.02e-06 ps=1.18554e-06 nrd=0.121951 nrs=0.219953 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=61940 $Y=41290 $D=28
M4982 216 4505 4506 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.12e-06 sb=1.95634e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=62260 $Y=41290 $D=28
M4983 4507 4505 216 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=1.6e-06 sb=1.47634e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=62740 $Y=41290 $D=28
M4984 VSS 162 4507 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=8.2e-14 pd=1.18e-06 ps=1.02e-06 nrd=0.219512 nrs=0.121951 sa=1.92e-06 sb=1.15634e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=63060 $Y=41290 $D=28
M4985 4508 162 VSS VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.2e-14 as=1.476e-13 pd=1.02e-06 ps=1.18e-06 nrd=0.121951 nrs=0.219512 sa=2e-06 sb=6.76341e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=63540 $Y=41290 $D=28
M4986 216 4505 4508 VSS lpnfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.922e-13 as=8.2e-14 pd=2.38e-06 ps=1.02e-06 nrd=0.434563 nrs=0.121951 sa=2e-06 sb=3.56341e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=63860 $Y=41290 $D=28
M4987 4510 4511 VSS VSS lpnfet w=8.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.602e-13 as=2.848e-13 pd=1.25e-06 ps=2.42e-06 nrd=0.202247 nrs=0.359551 sa=3.2e-07 sb=1.43191e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=20020 $Y=19590 $D=28
M4988 VSS 4511 4510 VSS lpnfet w=8.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87828e-13 as=1.602e-13 pd=1.40871e-06 ps=1.25e-06 nrd=0.237127 nrs=0.202247 sa=8e-07 sb=9.5191e-07 sd=0 panw1=0 panw2=3.9e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.49e-14 panw10=0 $X=20500 $Y=19590 $D=28
M4989 4509 106 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.144e-13 as=1.56172e-13 pd=2.6e-06 ps=1.17129e-06 nrd=0.756757 nrs=0.285193 sa=1.32e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.28e-14 panw10=0 $X=21020 $Y=19590 $D=28
M4990 4510 4509 126 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=2.752e-13 pd=1.22e-06 ps=2.36e-06 nrd=0.209302 nrs=0.372093 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=22200 $Y=19590 $D=28
M4991 126 4509 4510 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55095e-13 as=1.548e-13 pd=1.22857e-06 ps=1.22e-06 nrd=0.209701 nrs=0.209302 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=22680 $Y=19590 $D=28
M4992 4511 106 126 VSS lpnfet w=8.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.602e-13 as=1.60505e-13 pd=1.25e-06 ps=1.27143e-06 nrd=0.202247 nrs=0.202632 sa=1.2436e-06 sb=8e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=23160 $Y=19590 $D=28
M4993 126 106 4511 VSS lpnfet w=8.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.848e-13 as=1.602e-13 pd=2.42e-06 ps=1.25e-06 nrd=0.359551 nrs=0.202247 sa=1.7236e-06 sb=3.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=23640 $Y=19590 $D=28
M4994 4513 106 4512 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.8e-14 as=1.536e-13 pd=6.8e-07 ps=1.6e-06 nrd=0.208333 nrs=0.666667 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=24760 $Y=20000 $D=28
M4995 VSS 100 4513 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.92e-14 as=4.8e-14 pd=9.48148e-07 ps=6.8e-07 nrd=0.430556 nrs=0.208333 sa=6.4e-07 sb=1.72e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=25080 $Y=20000 $D=28
M4996 4511 100 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=1.77733e-13 pd=1.22e-06 ps=1.69877e-06 nrd=0.209302 nrs=0.24031 sa=7.15814e-07 sb=1.28e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.28e-14 panw10=0 $X=25520 $Y=19620 $D=28
M4997 VSS 100 4511 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=1.548e-13 pd=1.22e-06 ps=1.22e-06 nrd=0.209302 nrs=0.209302 sa=1.19581e-06 sb=8e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.28e-14 panw10=0 $X=26000 $Y=19620 $D=28
M4998 4511 100 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.752e-13 as=1.548e-13 pd=2.36e-06 ps=1.22e-06 nrd=0.372093 nrs=0.209302 sa=1.65349e-06 sb=3.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.28e-14 panw10=0 $X=26480 $Y=19620 $D=28
M4999 90 4512 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.944e-13 pd=2.48e-06 ps=2.48e-06 nrd=0.347826 nrs=0.347826 sa=3.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=27470 $Y=19590 $D=28
M5000 4515 4516 VSS VSS lpnfet w=8.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.602e-13 as=2.848e-13 pd=1.25e-06 ps=2.42e-06 nrd=0.202247 nrs=0.359551 sa=3.2e-07 sb=1.43191e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=52420 $Y=33990 $D=28
M5001 VSS 4516 4515 VSS lpnfet w=8.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87828e-13 as=1.602e-13 pd=1.40871e-06 ps=1.25e-06 nrd=0.237127 nrs=0.202247 sa=8e-07 sb=9.5191e-07 sd=0 panw1=0 panw2=3.9e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.49e-14 panw10=0 $X=52900 $Y=33990 $D=28
M5002 4514 224 VSS VSS lpnfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.144e-13 as=1.56172e-13 pd=2.6e-06 ps=1.17129e-06 nrd=0.756757 nrs=0.285193 sa=1.32e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.28e-14 panw10=0 $X=53420 $Y=33990 $D=28
M5003 4515 4514 150 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=2.752e-13 pd=1.22e-06 ps=2.36e-06 nrd=0.209302 nrs=0.372093 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=54600 $Y=33990 $D=28
M5004 150 4514 4515 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55095e-13 as=1.548e-13 pd=1.22857e-06 ps=1.22e-06 nrd=0.209701 nrs=0.209302 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=55080 $Y=33990 $D=28
M5005 4516 224 150 VSS lpnfet w=8.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.602e-13 as=1.60505e-13 pd=1.25e-06 ps=1.27143e-06 nrd=0.202247 nrs=0.202632 sa=1.2436e-06 sb=8e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=55560 $Y=33990 $D=28
M5006 150 224 4516 VSS lpnfet w=8.9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.848e-13 as=1.602e-13 pd=2.42e-06 ps=1.25e-06 nrd=0.359551 nrs=0.202247 sa=1.7236e-06 sb=3.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=56040 $Y=33990 $D=28
M5007 4518 224 4517 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.8e-14 as=1.536e-13 pd=6.8e-07 ps=1.6e-06 nrd=0.208333 nrs=0.666667 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=57160 $Y=34400 $D=28
M5008 VSS 159 4518 VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.92e-14 as=4.8e-14 pd=9.48148e-07 ps=6.8e-07 nrd=0.430556 nrs=0.208333 sa=6.4e-07 sb=1.72e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=57480 $Y=34400 $D=28
M5009 4516 159 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=1.77733e-13 pd=1.22e-06 ps=1.69877e-06 nrd=0.209302 nrs=0.24031 sa=7.15814e-07 sb=1.28e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.28e-14 panw10=0 $X=57920 $Y=34020 $D=28
M5010 VSS 159 4516 VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=1.548e-13 pd=1.22e-06 ps=1.22e-06 nrd=0.209302 nrs=0.209302 sa=1.19581e-06 sb=8e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.28e-14 panw10=0 $X=58400 $Y=34020 $D=28
M5011 4516 159 VSS VSS lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.752e-13 as=1.548e-13 pd=2.36e-06 ps=1.22e-06 nrd=0.372093 nrs=0.209302 sa=1.65349e-06 sb=3.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.28e-14 panw10=0 $X=58880 $Y=34020 $D=28
M5012 223 4517 VSS VSS lpnfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.944e-13 pd=2.48e-06 ps=2.48e-06 nrd=0.347826 nrs=0.347826 sa=3.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=59870 $Y=33990 $D=28
M5013 VSS 101 4519 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.63333e-14 as=9.44e-14 pd=8.2e-07 ps=1.28e-06 nrd=2.15833 nrs=2.36 sa=3.6e-07 sb=1.18e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=32160 $Y=32350 $D=28
M5014 4520 78 VSS VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4e-14 as=1.72667e-13 pd=6e-07 ps=1.64e-06 nrd=0.25 nrs=1.07917 sa=6.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=32700 $Y=32350 $D=28
M5015 102 4519 4520 VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28e-13 as=4e-14 pd=1.44e-06 ps=6e-07 nrd=0.8 nrs=0.25 sa=9.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=33020 $Y=32350 $D=28
M5016 VSS 217 4521 VSS lpnfet w=2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.63333e-14 as=9.44e-14 pd=8.2e-07 ps=1.28e-06 nrd=2.15833 nrs=2.36 sa=3.6e-07 sb=1.18e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=7.2e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=52560 $Y=25150 $D=28
M5017 4522 113 VSS VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4e-14 as=1.72667e-13 pd=6e-07 ps=1.64e-06 nrd=0.25 nrs=1.07917 sa=6.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=53100 $Y=25150 $D=28
M5018 814 4521 4522 VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.28e-13 as=4e-14 pd=1.44e-06 ps=6e-07 nrd=0.8 nrs=0.25 sa=9.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.92e-14 panw8=0 panw9=0 panw10=0 $X=53420 $Y=25150 $D=28
M5019 VSS data_in[0] 4523 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.06029e-13 as=9.6e-14 pd=8.85714e-07 ps=1.24e-06 nrd=1.1781 nrs=1.06667 sa=3.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=8910 $Y=18100 $D=28
M5020 101 4523 VSS VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.46e-14 as=1.66111e-13 pd=8.3e-07 ps=1.38762e-06 nrd=0.382979 nrs=0.751976 sa=6.89149e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=9470 $Y=17970 $D=28
M5021 VSS 4523 101 VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.18331e-13 as=8.46e-14 pd=1.8424e-06 ps=8.3e-07 nrd=0.988369 nrs=0.382979 sa=1.16915e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=9950 $Y=17970 $D=28
M5022 VSS weight_in[6] 4524 VSS lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.06029e-13 as=9.6e-14 pd=8.85714e-07 ps=1.24e-06 nrd=1.1781 nrs=1.06667 sa=3.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=1.2e-15 panw9=0 panw10=0 $X=46510 $Y=75700 $D=28
M5023 195 4524 VSS VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.46e-14 as=1.66111e-13 pd=8.3e-07 ps=1.38762e-06 nrd=0.382979 nrs=0.751976 sa=6.89149e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=47070 $Y=75570 $D=28
M5024 VSS 4524 195 VSS lpnfet w=4.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.18331e-13 as=8.46e-14 pd=1.8424e-06 ps=8.3e-07 nrd=0.988369 nrs=0.382979 sa=1.16915e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=47550 $Y=75570 $D=28
M5025 VSS data_in[7] 4525 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.198e-13 as=1.19e-13 pd=1.38e-06 ps=1.38e-06 nrd=1.03633 nrs=1.02941 sa=3.5e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=10840 $Y=56170 $D=28
M5026 186 4525 VSS VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.00696e-14 as=1.198e-13 pd=6.94783e-07 ps=1.38e-06 nrd=0.606138 nrs=1.03633 sa=7.9e-07 sb=8.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=11280 $Y=56170 $D=28
M5027 VSS 4525 186 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.61e-13 as=1.1953e-13 pd=2.08e-06 ps=1.18522e-06 nrd=0.775862 nrs=0.355322 sa=8.60345e-07 sb=3.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=9.6e-15 panw9=0 panw10=0 $X=11760 $Y=55930 $D=28
M5028 VSS weight_in[3] 4526 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.198e-13 as=1.19e-13 pd=1.38e-06 ps=1.38e-06 nrd=1.03633 nrs=1.02941 sa=3.5e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=34440 $Y=63370 $D=28
M5029 111 4526 VSS VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.00696e-14 as=1.198e-13 pd=6.94783e-07 ps=1.38e-06 nrd=0.606138 nrs=1.03633 sa=7.9e-07 sb=8.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=34880 $Y=63370 $D=28
M5030 VSS 4526 111 VSS lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.61e-13 as=1.1953e-13 pd=2.08e-06 ps=1.18522e-06 nrd=0.775862 nrs=0.355322 sa=8.60345e-07 sb=3.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=9.6e-15 panw9=0 panw10=0 $X=35360 $Y=63130 $D=28
M5031 945 37 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.44786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=3.36e-14 panw9=3.36e-14 panw10=0 $X=8860 $Y=73880 $D=111
M5032 872 874 945 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.12786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=9180 $Y=73880 $D=111
M5033 VDD 32 872 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.17896e-13 as=5.04e-14 pd=1.04901e-06 ps=6.4e-07 nrd=1.50377 nrs=0.642857 sa=1.17e-06 sb=6.47857e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=3.36e-14 $X=9660 $Y=73880 $D=111
M5034 VDD clk 870 VDD lppfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.18949e-13 as=1.664e-13 pd=1.94817e-06 ps=1.68e-06 nrd=0.809724 nrs=0.615385 sa=3.2e-07 sb=6.76154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=10180 $Y=74370 $D=111
M5035 VDD data_in[2] 871 VDD lppfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.51796e-13 as=1.98e-13 pd=1.07771e-06 ps=1.86e-06 nrd=0.421656 nrs=0.55 sa=3.3e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=10430 $Y=31090 $D=111
M5036 874 870 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.224e-13 as=1.43159e-13 pd=1.4e-06 ps=1.2738e-06 nrd=1.05882 nrs=1.2384 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=10690 $Y=74530 $D=111
M5037 141 871 VDD VDD lppfet w=9.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.746e-13 as=2.45404e-13 pd=1.33e-06 ps=1.74229e-06 nrd=0.185567 nrs=0.260818 sa=6.87835e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=10990 $Y=30720 $D=111
M5038 948 870 872 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.932e-13 pd=4.8e-07 ps=1.94e-06 nrd=0.357143 nrs=2.46429 sa=3.6e-07 sb=1.63357e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=11250 $Y=74050 $D=111
M5039 VDD 871 141 VDD lppfet w=9.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.104e-13 as=1.746e-13 pd=2.58e-06 ps=1.33e-06 nrd=0.329897 nrs=0.185567 sa=1.16784e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=11470 $Y=30720 $D=111
M5040 VDD 873 948 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.83789e-14 as=2.8e-14 pd=6.63158e-07 ps=4.8e-07 nrd=0.87218 nrs=0.357143 sa=6.8e-07 sb=1.41643e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=11570 $Y=74050 $D=111
M5041 873 872 VDD VDD lppfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.536e-13 as=1.17221e-13 pd=1.51e-06 ps=1.13684e-06 nrd=1.10069 nrs=0.508772 sa=8.53333e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=8.4e-15 panw8=2.4e-14 panw9=2.52e-14 panw10=0 $X=12110 $Y=73980 $D=111
M5042 875 870 873 VDD lppfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.74821e-13 as=2.536e-13 pd=1.37684e-06 ps=1.51e-06 nrd=0.758772 nrs=1.10069 sa=9.65625e-07 sb=1.3875e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.2e-14 panw10=1.56e-14 $X=12940 $Y=73660 $D=111
M5043 951 874 875 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=1.01979e-13 pd=4.9e-07 ps=8.03158e-07 nrd=0.375 nrs=1.30075 sa=1.70071e-06 sb=1.99036e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=13670 $Y=73860 $D=111
M5044 VDD 878 951 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.8e-14 as=2.94e-14 pd=6.22222e-07 ps=4.9e-07 nrd=1.25 nrs=0.375 sa=1.86714e-06 sb=1.67214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=14000 $Y=73860 $D=111
M5045 878 32 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=2.17e-13 pd=9.8e-07 ps=1.37778e-06 nrd=0.290323 nrs=0.564516 sa=1.19387e-06 sb=1.00097e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=4.8e-14 panw10=2.4e-14 $X=14730 $Y=73590 $D=111
M5046 VDD 875 878 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.49117e-13 as=1.116e-13 pd=1.53267e-06 ps=9.8e-07 nrd=0.648067 nrs=0.290323 sa=1.4571e-06 sb=5.20968e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=4.8e-14 panw10=2.4e-14 $X=15210 $Y=73590 $D=111
M5047 876 878 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=2.49117e-13 pd=1.88e-06 ps=1.53267e-06 nrd=0.516129 nrs=0.648067 sa=6.41129e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=7.2e-15 panw10=0 $X=15890 $Y=74130 $D=111
M5048 877 876 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=16830 $Y=73590 $D=111
M5049 VDD 876 877 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=17310 $Y=73590 $D=111
M5050 239 878 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=17790 $Y=73590 $D=111
M5051 VDD 878 239 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=18270 $Y=73590 $D=111
M5052 VDD clk 879 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.00267e-13 as=1.008e-13 pd=9.11111e-07 ps=1.28e-06 nrd=1.27891 nrs=1.28571 sa=3.6e-07 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=20160 $Y=17010 $D=111
M5053 954 clk VDD VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.04197e-13 as=2.50667e-13 pd=1.12459e-06 ps=2.27778e-06 nrd=0.212646 nrs=0.511565 sa=4.88571e-07 sb=5.86286e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=20640 $Y=16590 $D=111
M5054 882 884 954 VDD lppfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.664e-13 as=7.74033e-14 pd=1.68e-06 ps=8.3541e-07 nrd=0.615385 nrs=0.286255 sa=9.63077e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-15 panw9=0 panw10=0 $X=21040 $Y=16770 $D=111
M5055 880 95 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=8.05726e-14 pd=1.28e-06 ps=6.70502e-07 nrd=1.28571 nrs=1.02771 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=3.36e-14 panw8=0 panw9=0 panw10=0 $X=21850 $Y=16670 $D=111
M5056 VDD 879 884 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.41718e-13 as=2.688e-13 pd=2.01151e-06 ps=2.32e-06 nrd=0.34257 nrs=0.380952 sa=3.2e-07 sb=8.63095e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=22760 $Y=16310 $D=111
M5057 955 884 VDD VDD lppfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.2e-14 as=1.72656e-13 pd=8.4e-07 ps=1.43679e-06 nrd=0.2 nrs=0.479599 sa=7.58e-07 sb=7.68e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=23250 $Y=16250 $D=111
M5058 881 880 955 VDD lppfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.74273e-13 as=7.2e-14 pd=1.70455e-06 ps=8.4e-07 nrd=0.484091 nrs=0.2 sa=1.118e-06 sb=4.32e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=23610 $Y=16250 $D=111
M5059 957 882 881 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=8.13273e-14 pd=4.8e-07 ps=7.95455e-07 nrd=0.357143 nrs=1.03734 sa=4.57143e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=24140 $Y=16810 $D=111
M5060 VDD 883 957 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.67947e-14 as=2.8e-14 pd=7.60789e-07 ps=4.8e-07 nrd=0.851974 nrs=0.357143 sa=7.74286e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=24460 $Y=16810 $D=111
M5061 883 881 VDD VDD lppfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.64e-14 as=1.14505e-13 pd=8.4e-07 ps=1.30421e-06 nrd=0.375 nrs=0.496985 sa=7.71667e-07 sb=1.35583e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=24900 $Y=16610 $D=111
M5062 VDD 881 883 VDD lppfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.14505e-13 as=8.64e-14 pd=1.30421e-06 ps=8.4e-07 nrd=0.496985 nrs=0.375 sa=1.21167e-06 sb=8.75833e-07 sd=0 panw1=0 panw2=0 panw3=2.8e-15 panw4=3.5e-15 panw5=3.5e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.18e-14 panw9=0 panw10=0 $X=25380 $Y=16610 $D=111
M5063 883 68 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.832e-14 as=6.67947e-14 pd=6.16e-07 ps=7.60789e-07 nrd=0.871429 nrs=0.851974 sa=1.98286e-06 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=25870 $Y=16810 $D=111
M5064 887 882 883 VDD lppfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.2448e-13 pd=2.48e-06 ps=2.024e-06 nrd=0.347826 nrs=0.265217 sa=8.05217e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.64e-14 panw10=0 $X=26390 $Y=16370 $D=111
M5065 962 886 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.904e-13 pd=4.8e-07 ps=1.92e-06 nrd=0.357143 nrs=2.42857 sa=3.6e-07 sb=1.66286e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=9.6e-15 panw9=2.4e-14 panw10=0 $X=27430 $Y=16390 $D=111
M5066 887 884 962 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.16e-14 as=2.8e-14 pd=7.2e-07 ps=4.8e-07 nrd=0.785714 nrs=0.357143 sa=6.8e-07 sb=1.34286e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=9.6e-15 panw9=2.4e-14 panw10=0 $X=27750 $Y=16390 $D=111
M5067 VDD 68 887 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.792e-14 as=6.16e-14 pd=6.524e-07 ps=7.2e-07 nrd=1.12143 nrs=0.785714 sa=1.24e-06 sb=7.82857e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=9.6e-15 panw9=2.4e-14 panw10=0 $X=28310 $Y=16390 $D=111
M5068 VDD 887 886 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.792e-14 as=1.008e-13 pd=6.524e-07 ps=1.28e-06 nrd=1.12143 nrs=1.28571 sa=3.6e-07 sb=7.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=28630 $Y=17010 $D=111
M5069 100 887 VDD VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=2.3236e-13 pd=2.12e-06 ps=1.7242e-06 nrd=0.432432 nrs=0.424324 sa=7.18919e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=29070 $Y=16550 $D=111
M5070 889 888 VDD VDD lppfet w=9.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.746e-13 as=2.81222e-13 pd=1.33e-06 ps=2.99536e-06 nrd=0.185567 nrs=0.298887 sa=2.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=30330 $Y=71510 $D=111
M5071 VDD 105 889 VDD lppfet w=9.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.746e-13 as=1.746e-13 pd=1.33e-06 ps=1.33e-06 nrd=0.185567 nrs=0.185567 sa=7.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=30810 $Y=71510 $D=111
M5072 889 105 VDD VDD lppfet w=9.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.746e-13 as=1.746e-13 pd=1.33e-06 ps=1.33e-06 nrd=0.185567 nrs=0.185567 sa=1.2e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=31290 $Y=71510 $D=111
M5073 VDD 888 889 VDD lppfet w=9.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.10037e-13 as=1.746e-13 pd=1.44853e-06 ps=1.33e-06 nrd=0.22323 nrs=0.185567 sa=1.68e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=31770 $Y=71510 $D=111
M5074 402 889 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.77163e-13 pd=1.64e-06 ps=1.91147e-06 nrd=0.140625 nrs=0.169167 sa=1.59312e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=32290 $Y=71510 $D=111
M5075 VDD 889 402 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.70938e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=32770 $Y=71510 $D=111
M5076 402 889 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.82562e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=33250 $Y=71510 $D=111
M5077 VDD 889 402 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=1.94187e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=33730 $Y=71510 $D=111
M5078 190 890 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=1.34571e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=36480 $Y=66390 $D=111
M5079 VDD 807 190 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.835e-13 as=2.268e-13 pd=1.773e-06 ps=1.62e-06 nrd=0.178571 nrs=0.142857 sa=8.4e-07 sb=8.65714e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=36960 $Y=66390 $D=111
M5080 190 161 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.852e-13 as=2.835e-13 pd=3.16e-06 ps=1.773e-06 nrd=0.24263 nrs=0.178571 sa=1.4e-06 sb=3.05714e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=37520 $Y=66390 $D=111
M5081 891 147 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.15e-13 as=8.7e-14 pd=1.35e-06 ps=9.3913e-07 nrd=1.27778 nrs=0.966667 sa=2.6e-07 sb=1.62e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=38880 $Y=16930 $D=111
M5082 VDD 143 891 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.7e-14 as=1.15e-13 pd=9.3913e-07 ps=1.35e-06 nrd=0.966667 nrs=1.27778 sa=7.2e-07 sb=1.16e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=39340 $Y=16930 $D=111
M5083 125 154 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.664e-13 as=1.856e-13 pd=1.67e-06 ps=2.00348e-06 nrd=0.40625 nrs=0.453125 sa=6.9125e-07 sb=7e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=39800 $Y=16590 $D=111
M5084 892 153 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.16e-13 pd=1.66e-06 ps=3.24e-06 nrd=0.138462 nrs=0.246154 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=40010 $Y=73590 $D=111
M5085 VDD 891 125 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.35965e-13 as=1.664e-13 pd=2.62957e-06 ps=1.67e-06 nrd=0.576087 nrs=0.40625 sa=1.13125e-06 sb=2.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=40240 $Y=16590 $D=111
M5086 VDD 153 892 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=2.34e-13 pd=1.66e-06 ps=1.66e-06 nrd=0.138462 nrs=0.138462 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=40490 $Y=73590 $D=111
M5087 135 892 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=2.34e-13 pd=1.66e-06 ps=1.66e-06 nrd=0.138462 nrs=0.138462 sa=1.28e-06 sb=1.92246e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=40970 $Y=73590 $D=111
M5088 VDD 892 135 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=2.34e-13 pd=1.66e-06 ps=1.66e-06 nrd=0.138462 nrs=0.138462 sa=1.76e-06 sb=1.81908e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=41450 $Y=73590 $D=111
M5089 135 892 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=2.34e-13 pd=1.66e-06 ps=1.66e-06 nrd=0.138462 nrs=0.138462 sa=2e-06 sb=1.54308e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=41930 $Y=73590 $D=111
M5090 VDD 892 135 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37138e-13 as=2.34e-13 pd=1.86034e-06 ps=1.66e-06 nrd=0.140318 nrs=0.138462 sa=2e-06 sb=1.06308e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=42410 $Y=73590 $D=111
M5091 135 892 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.836e-13 as=1.86062e-13 pd=1.38e-06 ps=1.45966e-06 nrd=0.176471 nrs=0.178837 sa=2e-06 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.84e-14 panw10=0 $X=42890 $Y=73870 $D=111
M5092 VDD 892 135 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.468e-13 as=1.836e-13 pd=2.72e-06 ps=1.38e-06 nrd=0.333333 nrs=0.176471 sa=2e-06 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.84e-14 panw10=0 $X=43370 $Y=73870 $D=111
M5093 VDD 897 896 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.14842e-13 as=4.096e-13 pd=2.28299e-06 ps=3.2e-06 nrd=0.192164 nrs=0.25 sa=3.2e-07 sb=5.95469e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=60040 $Y=23190 $D=111
M5094 895 227 VDD VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.65e-13 as=1.22985e-13 pd=1.66e-06 ps=8.91791e-07 nrd=0.66 nrs=0.49194 sa=8.7e-07 sb=3.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.92e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=60590 $Y=23650 $D=111
M5095 244 227 896 VDD lppfet w=1.24e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.232e-13 as=3.968e-13 pd=1.6e-06 ps=3.12e-06 nrd=0.145161 nrs=0.258065 sa=3.2e-07 sb=1.82992e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=61540 $Y=23190 $D=111
M5096 897 895 244 VDD lppfet w=1.24e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.80872e-13 as=2.232e-13 pd=1.90929e-06 ps=1.6e-06 nrd=0.247705 nrs=0.145161 sa=8e-07 sb=1.49895e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=62020 $Y=23190 $D=111
M5097 VDD 264 897 VDD lppfet w=1.15e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.70201e-13 as=3.53228e-13 pd=1.97564e-06 ps=1.77071e-06 nrd=0.204311 nrs=0.267091 sa=1.52e-06 sb=9.96696e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=62740 $Y=23190 $D=111
M5098 901 195 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.46657e-13 pd=1.14e-06 ps=2.66377e-06 nrd=0.230769 nrs=0.405418 sa=2.4e-07 sb=1.93846e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=63170 $Y=45190 $D=111
M5099 898 264 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.86e-14 as=6.5788e-14 pd=7.7e-07 ps=4.81026e-07 nrd=0.875 nrs=0.839133 sa=2e-06 sb=1.29e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.68e-14 panw10=1.68e-14 $X=63300 $Y=23250 $D=111
M5100 897 264 VDD VDD lppfet w=6.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.48023e-13 pd=1.9e-06 ps=1.08231e-06 nrd=0.507937 nrs=0.372948 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=63300 $Y=23710 $D=111
M5101 VDD 195 901 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.6753e-13 as=1.404e-13 pd=1.60239e-06 ps=1.14e-06 nrd=0.275362 nrs=0.230769 sa=7.2e-07 sb=1.63333e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=63650 $Y=45190 $D=111
M5102 VDD 227 898 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09613e-13 as=6.86e-14 pd=8.75705e-07 ps=7.7e-07 nrd=1.39813 nrs=0.875 sa=2e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.68e-14 panw10=1.68e-14 $X=63910 $Y=23250 $D=111
M5103 900 901 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.638e-13 as=1.6753e-13 pd=1.2e-06 ps=1.60239e-06 nrd=0.269231 nrs=0.275362 sa=1.16e-06 sb=1.19333e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=64090 $Y=45190 $D=111
M5104 VDD 898 205 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50545e-13 as=1.904e-13 pd=2.00161e-06 ps=1.92e-06 nrd=0.611682 nrs=0.464844 sa=2.975e-07 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=64350 $Y=23850 $D=111
M5105 VDD 901 900 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.83944e-13 as=1.638e-13 pd=1.55322e-06 ps=1.2e-06 nrd=0.302341 nrs=0.269231 sa=1.7e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=64630 $Y=45190 $D=111
M5106 899 187 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.46212e-13 pd=1.88e-06 ps=1.23461e-06 nrd=0.516129 nrs=0.380365 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=65070 $Y=45350 $D=111
M5107 900 187 245 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=66030 $Y=45050 $D=111
M5108 903 906 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.25437e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=66210 $Y=64330 $D=111
M5109 245 187 900 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=66510 $Y=45050 $D=111
M5110 VDD 906 903 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.06605e-13 as=2.304e-13 pd=1.97457e-06 ps=1.64e-06 nrd=0.187137 nrs=0.140625 sa=8e-07 sb=7.74375e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=66690 $Y=64330 $D=111
M5111 901 899 245 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=66990 $Y=45050 $D=111
M5112 902 266 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.264e-13 as=2.44326e-13 pd=2.68e-06 ps=1.57349e-06 nrd=0.313725 nrs=0.234838 sa=1.36e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=67250 $Y=64330 $D=111
M5113 245 899 901 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=67470 $Y=45050 $D=111
M5114 903 266 250 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=4.064e-13 pd=1.63e-06 ps=3.18e-06 nrd=0.141732 nrs=0.251969 sa=3.2e-07 sb=1.71551e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=68190 $Y=64340 $D=111
M5115 250 266 903 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.60923e-13 as=2.286e-13 pd=1.68337e-06 ps=1.63e-06 nrd=0.161772 nrs=0.141732 sa=8e-07 sb=1.23551e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=68670 $Y=64340 $D=111
M5116 906 902 250 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.62977e-13 pd=1.64e-06 ps=1.69663e-06 nrd=0.140625 nrs=0.160509 sa=1.32211e-06 sb=7.0625e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=69200 $Y=64330 $D=111
M5117 250 902 906 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.896e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.176758 nrs=0.140625 sa=1.80211e-06 sb=2.2625e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=69680 $Y=64330 $D=111
M5118 905 266 VDD VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.75e-14 as=2.63077e-13 pd=8.9e-07 ps=2.41026e-06 nrd=0.39 nrs=1.05231 sa=2.496e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=70540 $Y=64360 $D=111
M5119 VDD 260 905 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.09141e-13 as=9.75e-14 pd=9.94949e-07 ps=8.9e-07 nrd=0.436566 nrs=0.39 sa=7.596e-07 sb=1.69e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=6e-15 panw9=0 panw10=0 $X=71050 $Y=64360 $D=111
M5120 906 260 VDD VDD lppfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.16e-13 as=2.61939e-13 pd=1.56e-06 ps=2.38788e-06 nrd=0.15 nrs=0.181902 sa=6.52e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=71460 $Y=64360 $D=111
M5121 VDD 260 906 VDD lppfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.16e-13 as=2.16e-13 pd=1.56e-06 ps=1.56e-06 nrd=0.15 nrs=0.15 sa=1.132e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=71940 $Y=64360 $D=111
M5122 906 260 VDD VDD lppfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.84e-13 as=2.16e-13 pd=3.04e-06 ps=1.56e-06 nrd=0.266667 nrs=0.15 sa=1.558e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=72420 $Y=64360 $D=111
M5123 276 905 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.096e-13 pd=3.2e-06 ps=3.2e-06 nrd=0.25 nrs=0.25 sa=3.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=73440 $Y=64310 $D=111
M5124 973 342 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3e-13 as=4.16e-13 pd=1.5e-06 ps=3.24e-06 nrd=0.0769231 nrs=0.246154 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=85360 $Y=73590 $D=111
M5125 353 323 973 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=1.3e-13 pd=1.66e-06 ps=1.5e-06 nrd=0.138462 nrs=0.0769231 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=85680 $Y=73590 $D=111
M5126 VDD 301 907 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.5965e-13 as=1.088e-13 pd=1.5e-06 ps=1.32e-06 nrd=1.38106 nrs=0.941176 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=86020 $Y=38550 $D=111
M5127 975 323 353 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3e-13 as=2.34e-13 pd=1.5e-06 ps=1.66e-06 nrd=0.0769231 nrs=0.138462 sa=1.12e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=86160 $Y=73590 $D=111
M5128 VDD 342 975 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=1.3e-13 pd=1.66e-06 ps=1.5e-06 nrd=0.138462 nrs=0.0769231 sa=1.44e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=86480 $Y=73590 $D=111
M5129 907 232 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.12e-14 as=1.5965e-13 pd=7e-07 ps=1.5e-06 nrd=0.529412 nrs=1.38106 sa=8.4e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=86540 $Y=38550 $D=111
M5130 976 342 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3e-13 as=2.34e-13 pd=1.5e-06 ps=1.66e-06 nrd=0.0769231 nrs=0.138462 sa=1.92e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=86960 $Y=73590 $D=111
M5131 908 314 907 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.224e-13 as=6.12e-14 pd=1.4e-06 ps=7e-07 nrd=1.05882 nrs=0.529412 sa=1.32e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=87020 $Y=38550 $D=111
M5132 413 908 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.024e-13 pd=1.92e-06 ps=9.6e-07 nrd=0.5 nrs=0.25 sa=5.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=7.68e-14 $X=87030 $Y=37640 $D=111
M5133 353 323 976 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=1.3e-13 pd=1.66e-06 ps=1.5e-06 nrd=0.138462 nrs=0.0769231 sa=2e-06 sb=1.908e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=87280 $Y=73590 $D=111
M5134 977 323 353 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3e-13 as=2.34e-13 pd=1.5e-06 ps=1.66e-06 nrd=0.0769231 nrs=0.138462 sa=2e-06 sb=1.428e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=87760 $Y=73590 $D=111
M5135 VDD 342 977 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=1.3e-13 pd=1.66e-06 ps=1.5e-06 nrd=0.138462 nrs=0.0769231 sa=2e-06 sb=1.108e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=88080 $Y=73590 $D=111
M5136 978 342 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3e-13 as=2.34e-13 pd=1.5e-06 ps=1.66e-06 nrd=0.0769231 nrs=0.138462 sa=2e-06 sb=6.28e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=88560 $Y=73590 $D=111
M5137 353 323 978 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.004e-13 as=1.3e-13 pd=3.24e-06 ps=1.5e-06 nrd=0.236923 nrs=0.0769231 sa=2e-06 sb=3.08e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=88880 $Y=73590 $D=111
M5138 382 375 VDD VDD lppfet w=1.21e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.178e-13 as=3.872e-13 pd=1.57e-06 ps=3.06e-06 nrd=0.14876 nrs=0.264463 sa=3.2e-07 sb=1.90975e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=102820 $Y=59190 $D=111
M5139 VDD 379 382 VDD lppfet w=1.21e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.178e-13 as=2.178e-13 pd=1.57e-06 ps=1.57e-06 nrd=0.14876 nrs=0.14876 sa=8e-07 sb=1.85818e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=103300 $Y=59190 $D=111
M5140 382 391 VDD VDD lppfet w=1.21e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.2e-13 as=2.178e-13 pd=2.44e-06 ps=1.57e-06 nrd=0.423468 nrs=0.14876 sa=1.28e-06 sb=1.80661e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=103780 $Y=59190 $D=111
M5141 VDD 375 382 VDD lppfet w=1.21e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.72474e-13 as=6.2e-13 pd=1.72089e-06 ps=2.44e-06 nrd=0.186103 nrs=0.423468 sa=1.80661e-06 sb=1.4e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=105000 $Y=59190 $D=111
M5142 382 379 VDD VDD lppfet w=1.21e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.178e-13 as=2.72474e-13 pd=1.57e-06 ps=1.72089e-06 nrd=0.14876 nrs=0.186103 sa=1.86678e-06 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=105560 $Y=59190 $D=111
M5143 VDD 391 382 VDD lppfet w=1.21e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.15136e-13 as=2.178e-13 pd=2.98846e-06 ps=1.57e-06 nrd=0.283543 nrs=0.14876 sa=1.91835e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=106040 $Y=59190 $D=111
M5144 985 401 417 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.276e-13 as=3.712e-13 pd=1.38e-06 ps=2.96e-06 nrd=0.0948276 nrs=0.275862 sa=3.2e-07 sb=1.84897e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=106180 $Y=71510 $D=111
M5145 VDD 392 985 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.16e-13 as=1.276e-13 pd=1.64e-06 ps=1.38e-06 nrd=0.160523 nrs=0.0948276 sa=6.6e-07 sb=1.81379e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=106520 $Y=71510 $D=111
M5146 986 392 VDD VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.392e-13 as=2.16e-13 pd=1.4e-06 ps=1.64e-06 nrd=0.103448 nrs=0.160523 sa=1.05103e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=107000 $Y=71630 $D=111
M5147 417 401 986 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.088e-13 as=1.392e-13 pd=1.52e-06 ps=1.4e-06 nrd=0.155172 nrs=0.103448 sa=1.41103e-06 sb=1.94e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=107360 $Y=71630 $D=111
M5148 987 401 417 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16e-13 as=2.088e-13 pd=1.36e-06 ps=1.52e-06 nrd=0.0862069 nrs=0.155172 sa=1.89103e-06 sb=1.46e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=107840 $Y=71630 $D=111
M5149 VDD 392 987 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.088e-13 as=1.16e-13 pd=1.52e-06 ps=1.36e-06 nrd=0.155172 nrs=0.0862069 sa=1.94207e-06 sb=1.14e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=108160 $Y=71630 $D=111
M5150 988 392 VDD VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16e-13 as=2.088e-13 pd=1.36e-06 ps=1.52e-06 nrd=0.0862069 nrs=0.155172 sa=1.99172e-06 sb=6.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=108640 $Y=71630 $D=111
M5151 417 401 988 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.944e-13 as=1.16e-13 pd=3e-06 ps=1.36e-06 nrd=0.293103 nrs=0.0862069 sa=2e-06 sb=3.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=108960 $Y=71630 $D=111
M5152 989 448 VDD VDD lppfet w=1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1e-13 as=3.2e-13 pd=1.2e-06 ps=2.64e-06 nrd=0.1 nrs=0.32 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=119400 $Y=57110 $D=111
M5153 911 433 989 VDD lppfet w=1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8e-13 as=1e-13 pd=1.36e-06 ps=1.2e-06 nrd=0.18 nrs=0.1 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=119720 $Y=57110 $D=111
M5154 990 433 911 VDD lppfet w=1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1e-13 as=1.8e-13 pd=1.2e-06 ps=1.36e-06 nrd=0.1 nrs=0.18 sa=1.12e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=120200 $Y=57110 $D=111
M5155 VDD 448 990 VDD lppfet w=1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.32281e-13 as=1e-13 pd=1.50877e-06 ps=1.2e-06 nrd=0.232281 nrs=0.1 sa=1.44e-06 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=120520 $Y=57110 $D=111
M5156 443 911 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.97319e-13 pd=1.64e-06 ps=1.93123e-06 nrd=0.140625 nrs=0.181469 sa=1.6325e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=121080 $Y=57110 $D=111
M5157 VDD 911 443 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.7375e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=121560 $Y=57110 $D=111
M5158 443 911 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=1.8425e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=122040 $Y=57110 $D=111
M5159 545 523 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=4.898e-13 pd=1.63e-06 ps=3.32e-06 nrd=0.141732 nrs=0.303677 sa=3.85669e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=134990 $Y=52010 $D=111
M5160 VDD 523 545 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.286e-13 pd=1.63e-06 ps=1.63e-06 nrd=0.141732 nrs=0.141732 sa=8.65669e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=135470 $Y=52010 $D=111
M5161 545 523 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.286e-13 pd=1.63e-06 ps=1.63e-06 nrd=0.141732 nrs=0.141732 sa=1.34567e-06 sb=1.77e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=135950 $Y=52010 $D=111
M5162 VDD 523 545 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.286e-13 pd=1.63e-06 ps=1.63e-06 nrd=0.141732 nrs=0.141732 sa=1.82567e-06 sb=1.29e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=136430 $Y=52010 $D=111
M5163 545 523 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.286e-13 pd=1.63e-06 ps=1.63e-06 nrd=0.141732 nrs=0.141732 sa=2e-06 sb=8.1e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=136910 $Y=52010 $D=111
M5164 VDD 523 545 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.191e-13 as=2.286e-13 pd=3.2e-06 ps=1.63e-06 nrd=0.259843 nrs=0.141732 sa=2e-06 sb=3.3e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=137390 $Y=52010 $D=111
M5165 915 608 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=8.96e-14 pd=6.4e-07 ps=1.2e-06 nrd=0.642857 nrs=1.14286 sa=3.2e-07 sb=1.34e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=1.56e-14 panw8=0 panw9=0 panw10=0 $X=139620 $Y=64460 $D=111
M5166 VDD 556 915 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.30435e-14 as=5.04e-14 pd=6.45217e-07 ps=6.4e-07 nrd=0.931677 nrs=0.642857 sa=8e-07 sb=8.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=1.56e-14 panw8=0 panw9=0 panw10=0 $X=140100 $Y=64460 $D=111
M5167 548 915 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.66957e-13 pd=1.92e-06 ps=1.47478e-06 nrd=0.5 nrs=0.407609 sa=7.775e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=140640 $Y=64310 $D=111
M5168 VDD 567 916 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.32971e-13 as=2.048e-13 pd=1.26136e-06 ps=1.92e-06 nrd=0.324636 nrs=0.5 sa=3.2e-07 sb=1.36375e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=141610 $Y=64310 $D=111
M5169 561 553 VDD VDD lppfet w=1.14e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.052e-13 as=2.36854e-13 pd=1.5e-06 ps=2.2468e-06 nrd=0.157895 nrs=0.182252 sa=4.74386e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=142050 $Y=64460 $D=111
M5170 VDD 854 561 VDD lppfet w=1.14e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.052e-13 as=2.052e-13 pd=1.5e-06 ps=1.5e-06 nrd=0.157895 nrs=0.157895 sa=9.54386e-07 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=142530 $Y=64460 $D=111
M5171 561 916 VDD VDD lppfet w=1.14e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.648e-13 as=2.052e-13 pd=2.92e-06 ps=1.5e-06 nrd=0.280702 nrs=0.157895 sa=1.43439e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=143010 $Y=64460 $D=111
M5172 996 778 917 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8e-14 as=2.56e-13 pd=1e-06 ps=2.24e-06 nrd=0.125 nrs=0.4 sa=3.2e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=0 $X=181680 $Y=42850 $D=111
M5173 997 757 996 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8e-14 as=8e-14 pd=1e-06 ps=1e-06 nrd=0.125 nrs=0.125 sa=6.4e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=0 $X=182000 $Y=42850 $D=111
M5174 VDD 759 997 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.97831e-13 as=8e-14 pd=1.36271e-06 ps=1e-06 nrd=0.30911 nrs=0.125 sa=9.6e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.88e-14 panw10=0 $X=182320 $Y=42850 $D=111
M5175 867 917 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=3.16529e-13 pd=3.2e-06 ps=2.18034e-06 nrd=0.25 nrs=0.193194 sa=1.0675e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=182880 $Y=42710 $D=111
M5176 772 716 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.56e-14 as=2.8224e-13 pd=7.8e-07 ps=2.304e-06 nrd=0.428571 nrs=1.6 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.56e-14 panw8=0 panw9=0 panw10=0 $X=183280 $Y=16860 $D=111
M5177 VDD 765 772 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=7.56e-14 pd=1.56e-06 ps=7.8e-07 nrd=0.857143 nrs=0.428571 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.56e-14 panw8=0 panw9=0 panw10=0 $X=183760 $Y=16860 $D=111
M5178 137 119 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=34920 $Y=21110 $D=111
M5179 270 820 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=68120 $Y=38250 $D=111
M5180 821 268 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=69320 $Y=74250 $D=111
M5181 387 366 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=100520 $Y=74250 $D=111
M5182 471 474 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=125720 $Y=28310 $D=111
M5183 465 476 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=125720 $Y=67050 $D=111
M5184 478 506 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=126520 $Y=35510 $D=111
M5185 484 477 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=126920 $Y=28310 $D=111
M5186 489 488 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=128520 $Y=38250 $D=111
M5187 486 505 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=130920 $Y=31050 $D=111
M5188 547 519 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=134920 $Y=38250 $D=111
M5189 531 530 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=136120 $Y=38250 $D=111
M5190 914 536 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=139320 $Y=31050 $D=111
M5191 550 554 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=142520 $Y=31050 $D=111
M5192 529 568 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=143720 $Y=28310 $D=111
M5193 565 557 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=144120 $Y=57110 $D=111
M5194 572 566 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=145320 $Y=57110 $D=111
M5195 603 614 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=153320 $Y=59850 $D=111
M5196 630 597 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=153720 $Y=42710 $D=111
M5197 601 624 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=154120 $Y=52650 $D=111
M5198 639 646 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=154920 $Y=42710 $D=111
M5199 619 616 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=155320 $Y=52650 $D=111
M5200 635 633 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=158120 $Y=52650 $D=111
M5201 642 666 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=160520 $Y=45450 $D=111
M5202 648 673 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=160920 $Y=57110 $D=111
M5203 670 652 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=162120 $Y=67050 $D=111
M5204 640 687 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=163320 $Y=59850 $D=111
M5205 675 683 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=165720 $Y=31050 $D=111
M5206 698 679 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=166520 $Y=59850 $D=111
M5207 862 692 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=169720 $Y=67050 $D=111
M5208 759 690 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=171720 $Y=42710 $D=111
M5209 720 731 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=173320 $Y=35510 $D=111
M5210 709 717 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=173720 $Y=31050 $D=111
M5211 677 686 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=174120 $Y=71510 $D=111
M5212 757 712 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=175320 $Y=42710 $D=111
M5213 750 726 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=176520 $Y=42710 $D=111
M5214 728 725 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=176520 $Y=57110 $D=111
M5215 730 636 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=178120 $Y=71510 $D=111
M5216 748 716 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=178520 $Y=21110 $D=111
M5217 765 733 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=182120 $Y=16650 $D=111
M5218 707 783 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=184120 $Y=71510 $D=111
M5219 773 736 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=184920 $Y=52650 $D=111
M5220 918 723 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=185720 $Y=28310 $D=111
M5221 776 785 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=186120 $Y=71510 $D=111
M5222 786 784 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=6.4e-14 panw10=1.28e-14 $X=187320 $Y=71510 $D=111
M5223 1705 417 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=112560 $Y=71510 $D=111
M5224 422 431 1705 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=112880 $Y=71510 $D=111
M5225 1706 430 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=116960 $Y=59650 $D=111
M5226 438 437 1706 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=117280 $Y=59650 $D=111
M5227 1707 456 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=120960 $Y=30850 $D=111
M5228 458 471 1707 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=121280 $Y=30850 $D=111
M5229 1708 458 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=124960 $Y=35510 $D=111
M5230 472 489 1708 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=125280 $Y=35510 $D=111
M5231 1709 492 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=129760 $Y=38050 $D=111
M5232 488 497 1709 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=130080 $Y=38050 $D=111
M5233 1710 528 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=130960 $Y=35510 $D=111
M5234 516 519 1710 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=131280 $Y=35510 $D=111
M5235 1711 522 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=132160 $Y=30850 $D=111
M5236 510 509 1711 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=132480 $Y=30850 $D=111
M5237 1712 505 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=135760 $Y=28310 $D=111
M5238 528 529 1712 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=136080 $Y=28310 $D=111
M5239 1713 559 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=136560 $Y=64310 $D=111
M5240 539 608 1713 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=136880 $Y=64310 $D=111
M5241 1714 556 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=140560 $Y=59650 $D=111
M5242 549 608 1714 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=140880 $Y=59650 $D=111
M5243 1715 597 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=148560 $Y=57110 $D=111
M5244 581 588 1715 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=148880 $Y=57110 $D=111
M5245 1716 626 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=156560 $Y=52450 $D=111
M5246 673 624 1716 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=156880 $Y=52450 $D=111
M5247 1717 632 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=160160 $Y=42710 $D=111
M5248 666 639 1717 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=160480 $Y=42710 $D=111
M5249 1718 617 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=168160 $Y=66850 $D=111
M5250 686 657 1718 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=168480 $Y=66850 $D=111
M5251 1719 726 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=169360 $Y=38050 $D=111
M5252 703 675 1719 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=169680 $Y=38050 $D=111
M5253 1720 863 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=172960 $Y=57110 $D=111
M5254 685 695 1720 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=173280 $Y=57110 $D=111
M5255 1721 703 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=174160 $Y=49910 $D=111
M5256 710 713 1721 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=174480 $Y=49910 $D=111
M5257 1722 686 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=176560 $Y=71510 $D=111
M5258 745 730 1722 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=176880 $Y=71510 $D=111
M5259 1723 731 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=177760 $Y=42710 $D=111
M5260 737 712 1723 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=178080 $Y=42710 $D=111
M5261 1724 652 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=179360 $Y=64310 $D=111
M5262 783 744 1724 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=179680 $Y=64310 $D=111
M5263 1725 759 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=185760 $Y=38050 $D=111
M5264 788 778 1725 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=186080 $Y=38050 $D=111
M5265 1726 783 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.176e-13 panw10=0 $X=187360 $Y=59650 $D=111
M5266 769 785 1726 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.44e-14 panw9=6.72e-14 panw10=0 $X=187680 $Y=59650 $D=111
M5267 13 63 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=14120 $Y=49910 $D=111
M5268 42 52 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=16520 $Y=30410 $D=111
M5269 48 43 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=17320 $Y=52010 $D=111
M5270 46 133 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=17720 $Y=21110 $D=111
M5271 60 58 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=20120 $Y=66410 $D=111
M5272 67 81 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=24520 $Y=73610 $D=111
M5273 888 885 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=29320 $Y=71510 $D=111
M5274 128 117 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=34920 $Y=13910 $D=111
M5275 145 893 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=41320 $Y=35510 $D=111
M5276 193 181 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=48920 $Y=57110 $D=111
M5277 208 815 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=56920 $Y=16010 $D=111
M5278 219 237 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=58920 $Y=37610 $D=111
M5279 222 230 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=62920 $Y=64310 $D=111
M5280 818 215 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=64120 $Y=59210 $D=111
M5281 262 249 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=68920 $Y=23210 $D=111
M5282 823 272 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=70520 $Y=73610 $D=111
M5283 336 284 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=78520 $Y=37610 $D=111
M5284 310 339 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=82920 $Y=13910 $D=111
M5285 317 363 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=85720 $Y=57110 $D=111
M5286 326 339 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=91320 $Y=13910 $D=111
M5287 339 345 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=91320 $Y=16010 $D=111
M5288 393 376 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=103320 $Y=73610 $D=111
M5289 416 380 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=107320 $Y=52010 $D=111
M5290 431 473 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=113320 $Y=73610 $D=111
M5291 429 417 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=115320 $Y=71510 $D=111
M5292 450 427 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=119720 $Y=30410 $D=111
M5293 469 458 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=123720 $Y=35510 $D=111
M5294 462 844 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=125320 $Y=64310 $D=111
M5295 515 509 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=127720 $Y=35510 $D=111
M5296 493 456 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=131320 $Y=42710 $D=111
M5297 524 497 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=131320 $Y=44810 $D=111
M5298 850 479 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=134120 $Y=13910 $D=111
M5299 564 850 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=140120 $Y=16010 $D=111
M5300 594 523 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=144920 $Y=49910 $D=111
M5301 575 586 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=145720 $Y=59210 $D=111
M5302 592 586 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=149320 $Y=52010 $D=111
M5303 599 607 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=152920 $Y=57110 $D=111
M5304 622 617 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=156120 $Y=57110 $D=111
M5305 651 655 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=163320 $Y=23210 $D=111
M5306 657 576 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=163320 $Y=66410 $D=111
M5307 760 658 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=164520 $Y=30410 $D=111
M5308 671 703 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=165720 $Y=42710 $D=111
M5309 689 860 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=169320 $Y=30410 $D=111
M5310 696 695 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=174520 $Y=66410 $D=111
M5311 747 734 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=179720 $Y=57110 $D=111
M5312 771 867 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=184520 $Y=37610 $D=111
M5313 756 918 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.752e-13 $X=186920 $Y=28310 $D=111
M5314 1728 298 1727 VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.6e-14 as=1.152e-13 pd=5.6e-07 ps=1.36e-06 nrd=0.277778 nrs=0.888889 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=74880 $Y=21110 $D=111
M5315 VDD 274 1728 VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10736e-13 as=3.6e-14 pd=8.352e-07 ps=5.6e-07 nrd=0.854444 nrs=0.277778 sa=6.4e-07 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=75200 $Y=21110 $D=111
M5316 825 1727 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.96864e-13 pd=1.92e-06 ps=1.4848e-06 nrd=0.5 nrs=0.480625 sa=9.08125e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=75840 $Y=21110 $D=111
M5317 1730 569 1729 VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.6e-14 as=1.152e-13 pd=5.6e-07 ps=1.36e-06 nrd=0.277778 nrs=0.888889 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=144880 $Y=24130 $D=111
M5318 VDD 568 1730 VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10736e-13 as=3.6e-14 pd=8.352e-07 ps=5.6e-07 nrd=0.854444 nrs=0.277778 sa=6.4e-07 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=145200 $Y=24130 $D=111
M5319 558 1729 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.96864e-13 pd=1.92e-06 ps=1.4848e-06 nrd=0.5 nrs=0.480625 sa=9.08125e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=145840 $Y=23850 $D=111
M5320 1732 765 1731 VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.6e-14 as=1.152e-13 pd=5.6e-07 ps=1.36e-06 nrd=0.277778 nrs=0.888889 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=4.32e-14 $X=186880 $Y=16930 $D=111
M5321 VDD 716 1732 VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.10736e-13 as=3.6e-14 pd=8.352e-07 ps=5.6e-07 nrd=0.854444 nrs=0.277778 sa=6.4e-07 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=4.32e-14 $X=187200 $Y=16930 $D=111
M5322 770 1731 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.96864e-13 pd=1.92e-06 ps=1.4848e-06 nrd=0.5 nrs=0.480625 sa=9.08125e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.68e-14 panw8=8.08e-14 panw9=0 panw10=0 $X=187840 $Y=16650 $D=111
M5323 VDD 129 1733 VDD lppfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.57609e-13 as=1.856e-13 pd=1.07174e-06 ps=1.8e-06 nrd=0.468516 nrs=0.551724 sa=3.2e-07 sb=1.38448e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=55780 $Y=31070 $D=111
M5324 209 170 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=3.42391e-13 pd=1.62e-06 ps=2.32826e-06 nrd=0.142857 nrs=0.215666 sa=5.99365e-07 sb=8.54444e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=56340 $Y=30390 $D=111
M5325 VDD 1733 209 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.718e-13 as=2.268e-13 pd=3.32e-06 ps=1.62e-06 nrd=0.297178 nrs=0.142857 sa=1.07937e-06 sb=3.74444e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=56820 $Y=30390 $D=111
M5326 VDD 246 1736 VDD lppfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.57609e-13 as=1.856e-13 pd=1.07174e-06 ps=1.8e-06 nrd=0.468516 nrs=0.551724 sa=3.2e-07 sb=1.38448e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=65780 $Y=57150 $D=111
M5327 247 241 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=3.42391e-13 pd=1.62e-06 ps=2.32826e-06 nrd=0.142857 nrs=0.215666 sa=5.99365e-07 sb=8.54444e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=66340 $Y=57150 $D=111
M5328 VDD 1736 247 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.718e-13 as=2.268e-13 pd=3.32e-06 ps=1.62e-06 nrd=0.297178 nrs=0.142857 sa=1.07937e-06 sb=3.74444e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=66820 $Y=57150 $D=111
M5329 VDD 742 1739 VDD lppfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.57609e-13 as=1.856e-13 pd=1.07174e-06 ps=1.8e-06 nrd=0.468516 nrs=0.551724 sa=3.2e-07 sb=1.38448e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=186180 $Y=52670 $D=111
M5330 869 788 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=3.42391e-13 pd=1.62e-06 ps=2.32826e-06 nrd=0.142857 nrs=0.215666 sa=5.99365e-07 sb=8.54444e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.752e-13 $X=186740 $Y=51990 $D=111
M5331 VDD 1739 869 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.718e-13 as=2.268e-13 pd=3.32e-06 ps=1.62e-06 nrd=0.297178 nrs=0.142857 sa=1.07937e-06 sb=3.74444e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.752e-13 $X=187220 $Y=51990 $D=111
M5332 VDD 55 1742 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20008e-13 as=1.984e-13 pd=1.01918e-06 ps=1.88e-06 nrd=0.312196 nrs=0.516129 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=14480 $Y=71700 $D=111
M5333 1743 23 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.62592e-13 pd=1.04e-06 ps=1.38082e-06 nrd=0.119048 nrs=0.230431 sa=6.6119e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=14960 $Y=71700 $D=111
M5334 37 1742 1743 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=9.8119e-07 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=15280 $Y=71700 $D=111
M5335 1744 1742 37 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.46119e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=15760 $Y=71700 $D=111
M5336 VDD 23 1744 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=1.78119e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=16080 $Y=71700 $D=111
M5337 VDD 101 1745 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20008e-13 as=1.984e-13 pd=1.01918e-06 ps=1.88e-06 nrd=0.312196 nrs=0.516129 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=26880 $Y=30880 $D=111
M5338 1746 199 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.62592e-13 pd=1.04e-06 ps=1.38082e-06 nrd=0.119048 nrs=0.230431 sa=6.6119e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=27360 $Y=30660 $D=111
M5339 52 1745 1746 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=9.8119e-07 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=27680 $Y=30660 $D=111
M5340 1747 1745 52 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.46119e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=28160 $Y=30660 $D=111
M5341 VDD 199 1747 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=1.78119e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=28480 $Y=30660 $D=111
M5342 VDD 129 1748 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20008e-13 as=1.984e-13 pd=1.01918e-06 ps=1.88e-06 nrd=0.312196 nrs=0.516129 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=37280 $Y=42900 $D=111
M5343 1749 82 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.62592e-13 pd=1.04e-06 ps=1.38082e-06 nrd=0.119048 nrs=0.230431 sa=6.6119e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=37760 $Y=42900 $D=111
M5344 140 1748 1749 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=9.8119e-07 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=38080 $Y=42900 $D=111
M5345 1750 1748 140 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.46119e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=38560 $Y=42900 $D=111
M5346 VDD 82 1750 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=1.78119e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=38880 $Y=42900 $D=111
M5347 VDD 394 1751 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20008e-13 as=1.984e-13 pd=1.01918e-06 ps=1.88e-06 nrd=0.312196 nrs=0.516129 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=100480 $Y=57300 $D=111
M5348 1752 437 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.62592e-13 pd=1.04e-06 ps=1.38082e-06 nrd=0.119048 nrs=0.230431 sa=6.6119e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=100960 $Y=57300 $D=111
M5349 369 1751 1752 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=9.8119e-07 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=101280 $Y=57300 $D=111
M5350 1753 1751 369 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.46119e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=101760 $Y=57300 $D=111
M5351 VDD 437 1753 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=1.78119e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=102080 $Y=57300 $D=111
M5352 VDD 913 1754 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20008e-13 as=1.984e-13 pd=1.01918e-06 ps=1.88e-06 nrd=0.312196 nrs=0.516129 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=140880 $Y=66880 $D=111
M5353 1755 561 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.62592e-13 pd=1.04e-06 ps=1.38082e-06 nrd=0.119048 nrs=0.230431 sa=6.6119e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=141360 $Y=66660 $D=111
M5354 552 1754 1755 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=9.8119e-07 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=141680 $Y=66660 $D=111
M5355 1756 1754 552 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.46119e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=142160 $Y=66660 $D=111
M5356 VDD 561 1756 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=1.78119e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=142480 $Y=66660 $D=111
M5357 VDD 868 1757 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20008e-13 as=1.984e-13 pd=1.01918e-06 ps=1.88e-06 nrd=0.312196 nrs=0.516129 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=186080 $Y=35700 $D=111
M5358 1758 771 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.62592e-13 pd=1.04e-06 ps=1.38082e-06 nrd=0.119048 nrs=0.230431 sa=6.6119e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=186560 $Y=35700 $D=111
M5359 781 1757 1758 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=9.8119e-07 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=1.008e-13 $X=186880 $Y=35700 $D=111
M5360 1759 1757 781 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.46119e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.404e-13 panw10=0 $X=187360 $Y=35700 $D=111
M5361 VDD 771 1759 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=1.78119e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.44e-14 panw9=9e-14 panw10=0 $X=187680 $Y=35700 $D=111
M5362 VDD 869 1760 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.20008e-13 as=1.984e-13 pd=1.01918e-06 ps=1.88e-06 nrd=0.312196 nrs=0.516129 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=186080 $Y=42900 $D=111
M5363 1761 779 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.62592e-13 pd=1.04e-06 ps=1.38082e-06 nrd=0.119048 nrs=0.230431 sa=6.6119e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=0 $X=186560 $Y=42900 $D=111
M5364 782 1760 1761 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=9.8119e-07 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.96e-14 panw10=1.008e-13 $X=186880 $Y=42900 $D=111
M5365 1762 1760 782 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.46119e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.404e-13 panw10=0 $X=187360 $Y=42900 $D=111
M5366 VDD 779 1762 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=8.4e-14 pd=2.32e-06 ps=1.04e-06 nrd=0.380952 nrs=0.119048 sa=1.78119e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.44e-14 panw9=9e-14 panw10=0 $X=187680 $Y=42900 $D=111
M5367 1763 21 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.792e-13 pd=9.2e-07 ps=1.76e-06 nrd=0.321429 nrs=0.571429 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=5.2e-14 panw8=4.64e-14 panw9=0 panw10=0 $X=8810 $Y=35510 $D=111
M5368 VDD 17 1763 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50477e-13 as=1.008e-13 pd=1.04172e-06 ps=9.2e-07 nrd=0.479839 nrs=0.321429 sa=8e-07 sb=8.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=6.72e-14 panw10=0 $X=9290 $Y=35510 $D=111
M5369 38 1763 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=3.49323e-13 pd=3.24e-06 ps=2.41828e-06 nrd=0.246154 nrs=0.2067 sa=7.80769e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-13 $X=9840 $Y=35510 $D=111
M5370 1765 825 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.792e-13 pd=9.2e-07 ps=1.76e-06 nrd=0.321429 nrs=0.571429 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=75210 $Y=23930 $D=111
M5371 VDD 281 1765 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50477e-13 as=1.008e-13 pd=1.04172e-06 ps=9.2e-07 nrd=0.479839 nrs=0.321429 sa=8e-07 sb=8.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=75690 $Y=23930 $D=111
M5372 826 1765 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=3.49323e-13 pd=3.24e-06 ps=2.41828e-06 nrd=0.246154 nrs=0.2067 sa=7.80769e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=76240 $Y=23190 $D=111
M5373 1767 525 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.792e-13 pd=9.2e-07 ps=1.76e-06 nrd=0.321429 nrs=0.571429 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=129210 $Y=45530 $D=111
M5374 VDD 517 1767 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50477e-13 as=1.008e-13 pd=1.04172e-06 ps=9.2e-07 nrd=0.479839 nrs=0.321429 sa=8e-07 sb=8.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=129690 $Y=45530 $D=111
M5375 498 1767 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=3.49323e-13 pd=3.24e-06 ps=2.41828e-06 nrd=0.246154 nrs=0.2067 sa=7.80769e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=130240 $Y=44790 $D=111
M5376 1769 501 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.792e-13 pd=9.2e-07 ps=1.76e-06 nrd=0.321429 nrs=0.571429 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=130810 $Y=28310 $D=111
M5377 VDD 504 1769 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50477e-13 as=1.008e-13 pd=1.04172e-06 ps=9.2e-07 nrd=0.479839 nrs=0.321429 sa=8e-07 sb=8.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=131290 $Y=28310 $D=111
M5378 507 1769 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=3.49323e-13 pd=3.24e-06 ps=2.41828e-06 nrd=0.246154 nrs=0.2067 sa=7.80769e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=131840 $Y=28310 $D=111
M5379 1771 558 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.792e-13 pd=9.2e-07 ps=1.76e-06 nrd=0.321429 nrs=0.571429 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=143610 $Y=31130 $D=111
M5380 VDD 554 1771 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50477e-13 as=1.008e-13 pd=1.04172e-06 ps=9.2e-07 nrd=0.479839 nrs=0.321429 sa=8e-07 sb=8.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=144090 $Y=31130 $D=111
M5381 573 1771 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=3.49323e-13 pd=3.24e-06 ps=2.41828e-06 nrd=0.246154 nrs=0.2067 sa=7.80769e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=144640 $Y=30390 $D=111
M5382 1773 642 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.792e-13 pd=9.2e-07 ps=1.76e-06 nrd=0.321429 nrs=0.571429 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=159210 $Y=49910 $D=111
M5383 VDD 633 1773 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50477e-13 as=1.008e-13 pd=1.04172e-06 ps=9.2e-07 nrd=0.479839 nrs=0.321429 sa=8e-07 sb=8.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=159690 $Y=49910 $D=111
M5384 634 1773 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=3.49323e-13 pd=3.24e-06 ps=2.41828e-06 nrd=0.246154 nrs=0.2067 sa=7.80769e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=160240 $Y=49910 $D=111
M5385 1775 625 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.792e-13 pd=9.2e-07 ps=1.76e-06 nrd=0.321429 nrs=0.571429 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=164410 $Y=45530 $D=111
M5386 VDD 660 1775 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50477e-13 as=1.008e-13 pd=1.04172e-06 ps=9.2e-07 nrd=0.479839 nrs=0.321429 sa=8e-07 sb=8.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=164890 $Y=45530 $D=111
M5387 663 1775 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=3.49323e-13 pd=3.24e-06 ps=2.41828e-06 nrd=0.246154 nrs=0.2067 sa=7.80769e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=165440 $Y=44790 $D=111
M5388 1777 677 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.792e-13 pd=9.2e-07 ps=1.76e-06 nrd=0.321429 nrs=0.571429 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=166010 $Y=67130 $D=111
M5389 VDD 692 1777 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50477e-13 as=1.008e-13 pd=1.04172e-06 ps=9.2e-07 nrd=0.479839 nrs=0.321429 sa=8e-07 sb=8.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=166490 $Y=67130 $D=111
M5390 672 1777 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=3.49323e-13 pd=3.24e-06 ps=2.41828e-06 nrd=0.246154 nrs=0.2067 sa=7.80769e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=167040 $Y=66390 $D=111
M5391 1779 684 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.792e-13 pd=9.2e-07 ps=1.76e-06 nrd=0.321429 nrs=0.571429 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=168010 $Y=64310 $D=111
M5392 VDD 679 1779 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50477e-13 as=1.008e-13 pd=1.04172e-06 ps=9.2e-07 nrd=0.479839 nrs=0.321429 sa=8e-07 sb=8.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=168490 $Y=64310 $D=111
M5393 861 1779 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=3.49323e-13 pd=3.24e-06 ps=2.41828e-06 nrd=0.246154 nrs=0.2067 sa=7.80769e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=169040 $Y=64310 $D=111
M5394 1781 707 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.792e-13 pd=9.2e-07 ps=1.76e-06 nrd=0.321429 nrs=0.571429 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=177210 $Y=64310 $D=111
M5395 VDD 736 1781 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50477e-13 as=1.008e-13 pd=1.04172e-06 ps=9.2e-07 nrd=0.479839 nrs=0.321429 sa=8e-07 sb=8.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=177690 $Y=64310 $D=111
M5396 738 1781 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=3.49323e-13 pd=3.24e-06 ps=2.41828e-06 nrd=0.246154 nrs=0.2067 sa=7.80769e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=178240 $Y=64310 $D=111
M5397 1783 778 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.792e-13 pd=9.2e-07 ps=1.76e-06 nrd=0.321429 nrs=0.571429 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=179210 $Y=42710 $D=111
M5398 VDD 757 1783 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50477e-13 as=1.008e-13 pd=1.04172e-06 ps=9.2e-07 nrd=0.479839 nrs=0.321429 sa=8e-07 sb=8.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=179690 $Y=42710 $D=111
M5399 749 1783 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=3.49323e-13 pd=3.24e-06 ps=2.41828e-06 nrd=0.246154 nrs=0.2067 sa=7.80769e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=180240 $Y=42710 $D=111
M5400 1785 770 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.792e-13 pd=9.2e-07 ps=1.76e-06 nrd=0.321429 nrs=0.571429 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=184810 $Y=16730 $D=111
M5401 VDD 772 1785 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50477e-13 as=1.008e-13 pd=1.04172e-06 ps=9.2e-07 nrd=0.479839 nrs=0.321429 sa=8e-07 sb=8.7e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=185290 $Y=16730 $D=111
M5402 774 1785 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=3.49323e-13 pd=3.24e-06 ps=2.41828e-06 nrd=0.246154 nrs=0.2067 sa=7.80769e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=185840 $Y=15990 $D=111
M5403 1787 44 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=18430 $Y=52330 $D=111
M5404 43 124 1787 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=18750 $Y=52330 $D=111
M5405 1788 124 43 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=19230 $Y=52330 $D=111
M5406 VDD 44 1788 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=19550 $Y=52330 $D=111
M5407 1789 80 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=21230 $Y=66730 $D=111
M5408 65 81 1789 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=21550 $Y=66730 $D=111
M5409 1790 81 65 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=22030 $Y=66730 $D=111
M5410 VDD 80 1790 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=22350 $Y=66730 $D=111
M5411 1791 98 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=42430 $Y=50030 $D=111
M5412 146 107 1791 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=42750 $Y=50030 $D=111
M5413 1792 107 146 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=43230 $Y=50030 $D=111
M5414 VDD 98 1792 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=43550 $Y=50030 $D=111
M5415 1793 82 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=44430 $Y=50030 $D=111
M5416 156 131 1793 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=44750 $Y=50030 $D=111
M5417 1794 131 156 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=45230 $Y=50030 $D=111
M5418 VDD 82 1794 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=45550 $Y=50030 $D=111
M5419 1795 243 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=66830 $Y=23530 $D=111
M5420 249 244 1795 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=67150 $Y=23530 $D=111
M5421 1796 244 249 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=67630 $Y=23530 $D=111
M5422 VDD 243 1796 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=67950 $Y=23530 $D=111
M5423 1797 409 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=105630 $Y=42830 $D=111
M5424 357 378 1797 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=105950 $Y=42830 $D=111
M5425 1798 378 357 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=106430 $Y=42830 $D=111
M5426 VDD 409 1798 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=106750 $Y=42830 $D=111
M5427 1799 439 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=115630 $Y=73930 $D=111
M5428 442 431 1799 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=115950 $Y=73930 $D=111
M5429 1800 431 442 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=116430 $Y=73930 $D=111
M5430 VDD 439 1800 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=116750 $Y=73930 $D=111
M5431 1801 845 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=126430 $Y=37930 $D=111
M5432 497 480 1801 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=126750 $Y=37930 $D=111
M5433 1802 480 497 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=127230 $Y=37930 $D=111
M5434 VDD 845 1802 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=127550 $Y=37930 $D=111
M5435 1803 485 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=128030 $Y=57230 $D=111
M5436 494 487 1803 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=128350 $Y=57230 $D=111
M5437 1804 487 494 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=128830 $Y=57230 $D=111
M5438 VDD 485 1804 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=129150 $Y=57230 $D=111
M5439 1805 493 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=132430 $Y=42830 $D=111
M5440 492 470 1805 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=132750 $Y=42830 $D=111
M5441 1806 470 492 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=133230 $Y=42830 $D=111
M5442 VDD 493 1806 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=133550 $Y=42830 $D=111
M5443 1807 491 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=133230 $Y=21230 $D=111
M5444 852 514 1807 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=133550 $Y=21230 $D=111
M5445 1808 514 852 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=134030 $Y=21230 $D=111
M5446 VDD 491 1808 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=134350 $Y=21230 $D=111
M5447 1809 500 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=137230 $Y=37930 $D=111
M5448 540 535 1809 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=137550 $Y=37930 $D=111
M5449 1810 535 540 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=138030 $Y=37930 $D=111
M5450 VDD 500 1810 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=138350 $Y=37930 $D=111
M5451 1811 512 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=139230 $Y=45130 $D=111
M5452 669 497 1811 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=139550 $Y=45130 $D=111
M5453 1812 497 669 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=140030 $Y=45130 $D=111
M5454 VDD 512 1812 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=140350 $Y=45130 $D=111
M5455 1813 575 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=145230 $Y=66730 $D=111
M5456 856 590 1813 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=145550 $Y=66730 $D=111
M5457 1814 590 856 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=146030 $Y=66730 $D=111
M5458 VDD 575 1814 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=146350 $Y=66730 $D=111
M5459 1815 575 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=156430 $Y=66730 $D=111
M5460 858 705 1815 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=156750 $Y=66730 $D=111
M5461 1816 705 858 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=157230 $Y=66730 $D=111
M5462 VDD 575 1816 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=157550 $Y=66730 $D=111
M5463 1817 648 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=162030 $Y=57230 $D=111
M5464 636 667 1817 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=162350 $Y=57230 $D=111
M5465 1818 667 636 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=162830 $Y=57230 $D=111
M5466 VDD 648 1818 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=163150 $Y=57230 $D=111
M5467 1819 575 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=165630 $Y=73930 $D=111
M5468 859 644 1819 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=165950 $Y=73930 $D=111
M5469 1820 644 859 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=166430 $Y=73930 $D=111
M5470 VDD 575 1820 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=166750 $Y=73930 $D=111
M5471 1821 693 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=180030 $Y=16330 $D=111
M5472 754 767 1821 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=180350 $Y=16330 $D=111
M5473 1822 767 754 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=180830 $Y=16330 $D=111
M5474 VDD 693 1822 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=181150 $Y=16330 $D=111
M5475 1823 681 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=181630 $Y=59530 $D=111
M5476 762 777 1823 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=181950 $Y=59530 $D=111
M5477 1824 777 762 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=182430 $Y=59530 $D=111
M5478 VDD 681 1824 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=182750 $Y=59530 $D=111
M5479 1825 681 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.36e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=184030 $Y=42830 $D=111
M5480 864 768 1825 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.04e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=184350 $Y=42830 $D=111
M5481 1826 768 864 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=5.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=184830 $Y=42830 $D=111
M5482 VDD 681 1826 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.50439e-13 as=8.4e-14 pd=2.70584e-06 ps=1.04e-06 nrd=0.35493 nrs=0.119048 sa=1.44e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=185150 $Y=42830 $D=111
M5483 VDD 15 1827 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.224e-13 panw10=0 $X=9280 $Y=21110 $D=111
M5484 1827 29 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-13 $X=9680 $Y=21110 $D=111
M5485 VDD 29 1827 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=10160 $Y=21110 $D=111
M5486 1827 15 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=10600 $Y=21110 $D=111
M5487 VDD 15 1827 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=11080 $Y=21110 $D=111
M5488 1827 29 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=11620 $Y=21010 $D=111
M5489 63 799 1827 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=12100 $Y=21110 $D=111
M5490 1827 799 63 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=12580 $Y=21110 $D=111
M5491 63 799 1827 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=13060 $Y=21110 $D=111
M5492 VDD 207 1831 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=52080 $Y=16430 $D=111
M5493 1831 235 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=52480 $Y=15990 $D=111
M5494 VDD 235 1831 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=52960 $Y=16310 $D=111
M5495 1831 207 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=53400 $Y=16040 $D=111
M5496 VDD 207 1831 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=53880 $Y=16040 $D=111
M5497 1831 235 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=54420 $Y=16310 $D=111
M5498 118 208 1831 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=54900 $Y=16170 $D=111
M5499 1831 208 118 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=55380 $Y=16170 $D=111
M5500 118 208 1831 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=55860 $Y=16170 $D=111
M5501 VDD 405 1835 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=108080 $Y=30830 $D=111
M5502 1835 445 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=108480 $Y=30390 $D=111
M5503 VDD 445 1835 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=108960 $Y=30710 $D=111
M5504 1835 405 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=109400 $Y=30440 $D=111
M5505 VDD 405 1835 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=109880 $Y=30440 $D=111
M5506 1835 445 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=110420 $Y=30710 $D=111
M5507 834 409 1835 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=110900 $Y=30570 $D=111
M5508 1835 409 834 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=111380 $Y=30570 $D=111
M5509 834 409 1835 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=111860 $Y=30570 $D=111
M5510 VDD 467 1839 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=120480 $Y=64310 $D=111
M5511 1839 460 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=120880 $Y=64310 $D=111
M5512 VDD 460 1839 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=121360 $Y=64310 $D=111
M5513 1839 467 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=121800 $Y=64310 $D=111
M5514 VDD 467 1839 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=122280 $Y=64310 $D=111
M5515 1839 460 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=122820 $Y=64210 $D=111
M5516 495 462 1839 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=123300 $Y=64310 $D=111
M5517 1839 462 495 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=123780 $Y=64310 $D=111
M5518 495 462 1839 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=124260 $Y=64310 $D=111
M5519 VDD 545 1843 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=121680 $Y=38030 $D=111
M5520 1843 488 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=122080 $Y=37590 $D=111
M5521 VDD 488 1843 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=122560 $Y=37910 $D=111
M5522 1843 545 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=123000 $Y=37640 $D=111
M5523 VDD 545 1843 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=123480 $Y=37640 $D=111
M5524 1843 488 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=124020 $Y=37910 $D=111
M5525 441 506 1843 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=124500 $Y=37770 $D=111
M5526 1843 506 441 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=124980 $Y=37770 $D=111
M5527 441 506 1843 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=125460 $Y=37770 $D=111
M5528 VDD 404 1847 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=121680 $Y=74030 $D=111
M5529 1847 490 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=122080 $Y=73590 $D=111
M5530 VDD 490 1847 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=122560 $Y=73910 $D=111
M5531 1847 404 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=123000 $Y=73640 $D=111
M5532 VDD 404 1847 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=123480 $Y=73640 $D=111
M5533 1847 490 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=124020 $Y=73910 $D=111
M5534 842 482 1847 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=124500 $Y=73770 $D=111
M5535 1847 482 842 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=124980 $Y=73770 $D=111
M5536 842 482 1847 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=125460 $Y=73770 $D=111
M5537 VDD 499 1851 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=124080 $Y=30830 $D=111
M5538 1851 472 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=124480 $Y=30390 $D=111
M5539 VDD 472 1851 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=124960 $Y=30710 $D=111
M5540 1851 499 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=125400 $Y=30440 $D=111
M5541 VDD 499 1851 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=125880 $Y=30440 $D=111
M5542 1851 472 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=126420 $Y=30710 $D=111
M5543 483 459 1851 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=126900 $Y=30570 $D=111
M5544 1851 459 483 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=127380 $Y=30570 $D=111
M5545 483 459 1851 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=127860 $Y=30570 $D=111
M5546 VDD 499 1855 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=132480 $Y=35510 $D=111
M5547 1855 516 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=132880 $Y=35510 $D=111
M5548 VDD 516 1855 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=133360 $Y=35510 $D=111
M5549 1855 499 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=133800 $Y=35510 $D=111
M5550 VDD 499 1855 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=134280 $Y=35510 $D=111
M5551 1855 516 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=134820 $Y=35410 $D=111
M5552 571 537 1855 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=135300 $Y=35510 $D=111
M5553 1855 537 571 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=135780 $Y=35510 $D=111
M5554 571 537 1855 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=136260 $Y=35510 $D=111
M5555 VDD 545 1859 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=139280 $Y=38030 $D=111
M5556 1859 547 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=139680 $Y=37590 $D=111
M5557 VDD 547 1859 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=140160 $Y=37910 $D=111
M5558 1859 545 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=140600 $Y=37640 $D=111
M5559 VDD 545 1859 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=141080 $Y=37640 $D=111
M5560 1859 547 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=141620 $Y=37910 $D=111
M5561 542 531 1859 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=142100 $Y=37770 $D=111
M5562 1859 531 542 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=142580 $Y=37770 $D=111
M5563 542 531 1859 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=143060 $Y=37770 $D=111
M5564 VDD 545 1863 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=139280 $Y=57110 $D=111
M5565 1863 565 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=139680 $Y=57110 $D=111
M5566 VDD 565 1863 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=140160 $Y=57110 $D=111
M5567 1863 545 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=140600 $Y=57110 $D=111
M5568 VDD 545 1863 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=141080 $Y=57110 $D=111
M5569 1863 565 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=141620 $Y=57010 $D=111
M5570 583 572 1863 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=142100 $Y=57110 $D=111
M5571 1863 572 583 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=142580 $Y=57110 $D=111
M5572 583 572 1863 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=143060 $Y=57110 $D=111
M5573 VDD 562 1867 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=169280 $Y=49910 $D=111
M5574 1867 691 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=169680 $Y=49910 $D=111
M5575 VDD 691 1867 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=170160 $Y=49910 $D=111
M5576 1867 562 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=170600 $Y=49910 $D=111
M5577 VDD 562 1867 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=171080 $Y=49910 $D=111
M5578 1867 691 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=171620 $Y=49810 $D=111
M5579 702 739 1867 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=172100 $Y=49910 $D=111
M5580 1867 739 702 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=172580 $Y=49910 $D=111
M5581 702 739 1867 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=173060 $Y=49910 $D=111
M5582 VDD 742 1871 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=176480 $Y=30830 $D=111
M5583 1871 737 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=176880 $Y=30390 $D=111
M5584 VDD 737 1871 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=177360 $Y=30710 $D=111
M5585 1871 742 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=177800 $Y=30440 $D=111
M5586 VDD 742 1871 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=178280 $Y=30440 $D=111
M5587 1871 737 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=178820 $Y=30710 $D=111
M5588 764 741 1871 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=179300 $Y=30570 $D=111
M5589 1871 741 764 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=179780 $Y=30570 $D=111
M5590 764 741 1871 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=180260 $Y=30570 $D=111
M5591 VDD 729 1875 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=176880 $Y=59630 $D=111
M5592 1875 776 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=177280 $Y=59190 $D=111
M5593 VDD 776 1875 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=177760 $Y=59510 $D=111
M5594 1875 729 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=178200 $Y=59240 $D=111
M5595 VDD 729 1875 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=178680 $Y=59240 $D=111
M5596 1875 776 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=179220 $Y=59510 $D=111
M5597 751 786 1875 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=179700 $Y=59370 $D=111
M5598 1875 786 751 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=180180 $Y=59370 $D=111
M5599 751 786 1875 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=180660 $Y=59370 $D=111
M5600 VDD 729 1879 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=179280 $Y=71510 $D=111
M5601 1879 745 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=179680 $Y=71510 $D=111
M5602 VDD 745 1879 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=180160 $Y=71510 $D=111
M5603 1879 729 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=180600 $Y=71510 $D=111
M5604 VDD 729 1879 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=181080 $Y=71510 $D=111
M5605 1879 745 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=181620 $Y=71410 $D=111
M5606 763 758 1879 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=182100 $Y=71510 $D=111
M5607 1879 758 763 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=182580 $Y=71510 $D=111
M5608 763 758 1879 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-15 $X=183060 $Y=71510 $D=111
M5609 VDD 755 1883 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45582e-13 as=3.01e-13 pd=1.35464e-06 ps=2.42e-06 nrd=0.196838 nrs=0.406977 sa=3.5e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=184080 $Y=23630 $D=111
M5610 1883 742 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.37649e-13 as=2.20065e-13 pd=1.89298e-06 ps=2.04771e-06 nrd=0.140621 nrs=0.130216 sa=6.15538e-07 sb=1.55692e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=184480 $Y=23190 $D=111
M5611 VDD 742 1883 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80851e-13 as=1.79151e-13 pd=1.56956e-06 ps=1.42702e-06 nrd=0.188308 nrs=0.186538 sa=1.16265e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=184960 $Y=23510 $D=111
M5612 1883 755 VDD VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.25e-13 as=2.30677e-13 pd=1.61e-06 ps=2.00199e-06 nrd=0.144 nrs=0.147633 sa=1.30832e-06 sb=1.74512e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-14 $X=185400 $Y=23240 $D=111
M5613 VDD 755 1883 VDD lppfet w=1.25e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.97989e-13 as=2.25e-13 pd=2.02107e-06 ps=1.61e-06 nrd=0.190713 nrs=0.144 sa=1.68512e-06 sb=1.64144e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=185880 $Y=23240 $D=111
M5614 1883 742 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.02255e-13 as=2.57462e-13 pd=1.55127e-06 ps=1.74621e-06 nrd=0.173401 nrs=0.220732 sa=1.84259e-06 sb=1.61556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=186420 $Y=23510 $D=111
M5615 787 780 1883 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.09745e-13 pd=1.48e-06 ps=1.60873e-06 nrd=0.160714 nrs=0.167208 sa=1.785e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.488e-13 $X=186900 $Y=23370 $D=111
M5616 1883 780 787 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=2.016e-13 pd=1.48e-06 ps=1.48e-06 nrd=0.160714 nrs=0.160714 sa=1.845e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.824e-13 panw10=2.4e-15 $X=187380 $Y=23370 $D=111
M5617 787 780 1883 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=2.016e-13 pd=2.88e-06 ps=1.48e-06 nrd=0.285714 nrs=0.160714 sa=1.905e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=6.88e-14 panw8=1.136e-13 panw9=4.8e-14 panw10=2.4e-15 $X=187860 $Y=23370 $D=111
M5618 VDD 411 1887 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=104670 $Y=74030 $D=111
M5619 1887 387 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=105150 $Y=74030 $D=111
M5620 VDD 387 1887 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.28e-06 sb=1.76e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=105630 $Y=74030 $D=111
M5621 1887 411 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.76e-06 sb=1.28e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=106110 $Y=74030 $D=111
M5622 383 393 1887 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=106590 $Y=74030 $D=111
M5623 1887 393 383 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=107070 $Y=74030 $D=111
M5624 VDD 422 1890 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=108670 $Y=64330 $D=111
M5625 1890 411 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=109150 $Y=64330 $D=111
M5626 VDD 411 1890 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.28e-06 sb=1.76e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=109630 $Y=64330 $D=111
M5627 1890 422 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.76e-06 sb=1.28e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=110110 $Y=64330 $D=111
M5628 833 420 1890 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=110590 $Y=64330 $D=111
M5629 1890 420 833 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=111070 $Y=64330 $D=111
M5630 VDD 411 1893 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=117870 $Y=74030 $D=111
M5631 1893 442 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=118350 $Y=74030 $D=111
M5632 VDD 442 1893 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.28e-06 sb=1.76e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=118830 $Y=74030 $D=111
M5633 1893 411 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.76e-06 sb=1.28e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=119310 $Y=74030 $D=111
M5634 464 840 1893 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=119790 $Y=74030 $D=111
M5635 1893 840 464 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=120270 $Y=74030 $D=111
M5636 VDD 518 1896 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=133470 $Y=57130 $D=111
M5637 1896 524 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=133950 $Y=57130 $D=111
M5638 VDD 524 1896 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.28e-06 sb=1.76e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=134430 $Y=57130 $D=111
M5639 1896 518 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.76e-06 sb=1.28e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=134910 $Y=57130 $D=111
M5640 511 534 1896 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=135390 $Y=57130 $D=111
M5641 1896 534 511 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=135870 $Y=57130 $D=111
M5642 VDD 912 1899 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=137070 $Y=42730 $D=111
M5643 1899 510 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=137550 $Y=42730 $D=111
M5644 VDD 510 1899 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.28e-06 sb=1.76e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=138030 $Y=42730 $D=111
M5645 1899 912 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.76e-06 sb=1.28e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=138510 $Y=42730 $D=111
M5646 532 546 1899 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=138990 $Y=42730 $D=111
M5647 1899 546 532 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=139470 $Y=42730 $D=111
M5648 VDD 594 1902 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=150270 $Y=49930 $D=111
M5649 1902 669 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=150750 $Y=49930 $D=111
M5650 VDD 669 1902 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.28e-06 sb=1.76e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=151230 $Y=49930 $D=111
M5651 1902 594 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.76e-06 sb=1.28e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=151710 $Y=49930 $D=111
M5652 587 598 1902 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=152190 $Y=49930 $D=111
M5653 1902 598 587 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=152670 $Y=49930 $D=111
M5654 VDD 562 1905 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=158670 $Y=66830 $D=111
M5655 1905 636 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=159150 $Y=66830 $D=111
M5656 VDD 636 1905 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.28e-06 sb=1.76e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=159630 $Y=66830 $D=111
M5657 1905 562 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.76e-06 sb=1.28e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=160110 $Y=66830 $D=111
M5658 857 674 1905 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=160590 $Y=66830 $D=111
M5659 1905 674 857 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=161070 $Y=66830 $D=111
M5660 VDD 518 1908 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=159470 $Y=52430 $D=111
M5661 1908 653 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=159950 $Y=52430 $D=111
M5662 VDD 653 1908 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.28e-06 sb=1.76e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=160430 $Y=52430 $D=111
M5663 1908 518 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.76e-06 sb=1.28e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=160910 $Y=52430 $D=111
M5664 637 650 1908 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=161390 $Y=52430 $D=111
M5665 1908 650 637 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=161870 $Y=52430 $D=111
M5666 VDD 598 1911 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=165870 $Y=49930 $D=111
M5667 1911 710 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=166350 $Y=49930 $D=111
M5668 VDD 710 1911 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.28e-06 sb=1.76e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=166830 $Y=49930 $D=111
M5669 1911 598 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.76e-06 sb=1.28e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=167310 $Y=49930 $D=111
M5670 690 727 1911 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=167790 $Y=49930 $D=111
M5671 1911 727 690 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=168270 $Y=49930 $D=111
M5672 VDD 674 1914 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=167870 $Y=59630 $D=111
M5673 1914 696 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=168350 $Y=59630 $D=111
M5674 VDD 696 1914 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.28e-06 sb=1.76e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=168830 $Y=59630 $D=111
M5675 1914 674 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.76e-06 sb=1.28e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=169310 $Y=59630 $D=111
M5676 784 728 1914 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=169790 $Y=59630 $D=111
M5677 1914 728 784 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=170270 $Y=59630 $D=111
M5678 VDD 518 1917 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=183870 $Y=59630 $D=111
M5679 1917 769 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=184350 $Y=59630 $D=111
M5680 VDD 769 1917 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.28e-06 sb=1.76e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=184830 $Y=59630 $D=111
M5681 1917 518 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=1.76e-06 sb=1.28e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=185310 $Y=59630 $D=111
M5682 866 775 1917 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=185790 $Y=59630 $D=111
M5683 1917 775 866 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=186270 $Y=59630 $D=111
M5684 1921 173 1920 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=2.544e-13 pd=8.6e-07 ps=2.16e-06 nrd=0.151515 nrs=0.584022 sa=3.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=47280 $Y=23830 $D=111
M5685 VDD 140 1921 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.07458e-13 as=6.6e-14 pd=1.22474e-06 ps=8.6e-07 nrd=0.476257 nrs=0.151515 sa=6.8e-07 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=47600 $Y=23830 $D=111
M5686 147 1920 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.02342e-13 pd=3.2e-06 ps=2.37526e-06 nrd=0.25 nrs=0.24557 sa=8.88906e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=48240 $Y=23210 $D=111
M5687 1923 486 1922 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=2.544e-13 pd=8.6e-07 ps=2.16e-06 nrd=0.151515 nrs=0.584022 sa=3.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=123280 $Y=23830 $D=111
M5688 VDD 474 1923 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.07458e-13 as=6.6e-14 pd=1.22474e-06 ps=8.6e-07 nrd=0.476257 nrs=0.151515 sa=6.8e-07 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=123600 $Y=23830 $D=111
M5689 501 1922 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.02342e-13 pd=3.2e-06 ps=2.37526e-06 nrd=0.25 nrs=0.24557 sa=8.88906e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=124240 $Y=23210 $D=111
M5690 1925 582 1924 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=2.544e-13 pd=8.6e-07 ps=2.16e-06 nrd=0.151515 nrs=0.584022 sa=3.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=147680 $Y=31030 $D=111
M5691 VDD 573 1925 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.07458e-13 as=6.6e-14 pd=1.22474e-06 ps=8.6e-07 nrd=0.476257 nrs=0.151515 sa=6.8e-07 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=148000 $Y=31030 $D=111
M5692 591 1924 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.02342e-13 pd=3.2e-06 ps=2.37526e-06 nrd=0.25 nrs=0.24557 sa=8.88906e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=148640 $Y=30410 $D=111
M5693 1927 622 1926 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=2.544e-13 pd=8.6e-07 ps=2.16e-06 nrd=0.151515 nrs=0.584022 sa=3.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=154480 $Y=64310 $D=111
M5694 VDD 609 1927 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.07458e-13 as=6.6e-14 pd=1.22474e-06 ps=8.6e-07 nrd=0.476257 nrs=0.151515 sa=6.8e-07 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=154800 $Y=64310 $D=111
M5695 602 1926 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.02342e-13 pd=3.2e-06 ps=2.37526e-06 nrd=0.25 nrs=0.24557 sa=8.88906e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=155440 $Y=64310 $D=111
M5696 1929 592 1928 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=2.544e-13 pd=8.6e-07 ps=2.16e-06 nrd=0.151515 nrs=0.584022 sa=3.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=155680 $Y=49910 $D=111
M5697 VDD 634 1929 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.07458e-13 as=6.6e-14 pd=1.22474e-06 ps=8.6e-07 nrd=0.476257 nrs=0.151515 sa=6.8e-07 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=156000 $Y=49910 $D=111
M5698 600 1928 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.02342e-13 pd=3.2e-06 ps=2.37526e-06 nrd=0.25 nrs=0.24557 sa=8.88906e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=156640 $Y=49910 $D=111
M5699 1931 592 1930 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=2.544e-13 pd=8.6e-07 ps=2.16e-06 nrd=0.151515 nrs=0.584022 sa=3.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=157680 $Y=38230 $D=111
M5700 VDD 663 1931 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.07458e-13 as=6.6e-14 pd=1.22474e-06 ps=8.6e-07 nrd=0.476257 nrs=0.151515 sa=6.8e-07 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=158000 $Y=38230 $D=111
M5701 574 1930 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.02342e-13 pd=3.2e-06 ps=2.37526e-06 nrd=0.25 nrs=0.24557 sa=8.88906e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=158640 $Y=37610 $D=111
M5702 1933 630 1932 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=2.544e-13 pd=8.6e-07 ps=2.16e-06 nrd=0.151515 nrs=0.584022 sa=3.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=158080 $Y=42710 $D=111
M5703 VDD 646 1933 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.07458e-13 as=6.6e-14 pd=1.22474e-06 ps=8.6e-07 nrd=0.476257 nrs=0.151515 sa=6.8e-07 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=158400 $Y=42710 $D=111
M5704 625 1932 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.02342e-13 pd=3.2e-06 ps=2.37526e-06 nrd=0.25 nrs=0.24557 sa=8.88906e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=159040 $Y=42710 $D=111
M5705 1935 670 1934 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=2.544e-13 pd=8.6e-07 ps=2.16e-06 nrd=0.151515 nrs=0.584022 sa=3.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=164480 $Y=59830 $D=111
M5706 VDD 576 1935 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.07458e-13 as=6.6e-14 pd=1.22474e-06 ps=8.6e-07 nrd=0.476257 nrs=0.151515 sa=6.8e-07 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=164800 $Y=59830 $D=111
M5707 684 1934 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.02342e-13 pd=3.2e-06 ps=2.37526e-06 nrd=0.25 nrs=0.24557 sa=8.88906e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=165440 $Y=59210 $D=111
M5708 1937 748 1936 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=2.544e-13 pd=8.6e-07 ps=2.16e-06 nrd=0.151515 nrs=0.584022 sa=3.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=182080 $Y=23830 $D=111
M5709 VDD 717 1937 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.07458e-13 as=6.6e-14 pd=1.22474e-06 ps=8.6e-07 nrd=0.476257 nrs=0.151515 sa=6.8e-07 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=182400 $Y=23830 $D=111
M5710 761 1936 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.02342e-13 pd=3.2e-06 ps=2.37526e-06 nrd=0.25 nrs=0.24557 sa=8.88906e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=183040 $Y=23210 $D=111
M5711 1939 750 1938 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.6e-14 as=2.544e-13 pd=8.6e-07 ps=2.16e-06 nrd=0.151515 nrs=0.584022 sa=3.6e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=182880 $Y=52630 $D=111
M5712 VDD 746 1939 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.07458e-13 as=6.6e-14 pd=1.22474e-06 ps=8.6e-07 nrd=0.476257 nrs=0.151515 sa=6.8e-07 sb=9.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=183200 $Y=52630 $D=111
M5713 732 1938 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.02342e-13 pd=3.2e-06 ps=2.37526e-06 nrd=0.25 nrs=0.24557 sa=8.88906e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=183840 $Y=52010 $D=111
M5714 34 52 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=12480 $Y=35510 $D=111
M5715 VDD 70 34 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=12960 $Y=35510 $D=111
M5716 19 40 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=14480 $Y=16650 $D=111
M5717 VDD 29 19 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=14960 $Y=16650 $D=111
M5718 35 30 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=15280 $Y=49910 $D=111
M5719 VDD 14 35 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=15760 $Y=49910 $D=111
M5720 31 36 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=16080 $Y=57110 $D=111
M5721 VDD 48 31 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=16560 $Y=57110 $D=111
M5722 36 44 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=17680 $Y=57110 $D=111
M5723 VDD 124 36 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=18160 $Y=57110 $D=111
M5724 61 44 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=20480 $Y=49910 $D=111
M5725 VDD 124 61 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=20960 $Y=49910 $D=111
M5726 64 91 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=20880 $Y=74250 $D=111
M5727 VDD 67 64 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=21360 $Y=74250 $D=111
M5728 116 132 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=37280 $Y=16650 $D=111
M5729 VDD 137 116 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=37760 $Y=16650 $D=111
M5730 154 140 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=45680 $Y=23850 $D=111
M5731 VDD 173 154 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=46160 $Y=23850 $D=111
M5732 243 198 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=54480 $Y=21110 $D=111
M5733 VDD 814 243 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=54960 $Y=21110 $D=111
M5734 816 815 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=58080 $Y=16650 $D=111
M5735 VDD 207 816 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=58560 $Y=16650 $D=111
M5736 258 243 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=65280 $Y=23850 $D=111
M5737 VDD 244 258 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=65760 $Y=23850 $D=111
M5738 259 258 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=70080 $Y=23850 $D=111
M5739 VDD 262 259 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=70560 $Y=23850 $D=111
M5740 277 904 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=70480 $Y=71510 $D=111
M5741 VDD 289 277 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=70960 $Y=71510 $D=111
M5742 281 274 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=73280 $Y=21110 $D=111
M5743 VDD 298 281 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=73760 $Y=21110 $D=111
M5744 292 297 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=76880 $Y=42710 $D=111
M5745 VDD 286 292 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=77360 $Y=42710 $D=111
M5746 909 361 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=96480 $Y=71510 $D=111
M5747 VDD 830 909 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=96960 $Y=71510 $D=111
M5748 391 363 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=96880 $Y=57110 $D=111
M5749 VDD 359 391 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=97360 $Y=57110 $D=111
M5750 372 376 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=101680 $Y=74250 $D=111
M5751 VDD 387 372 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=102160 $Y=74250 $D=111
M5752 414 438 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=107280 $Y=59850 $D=111
M5753 VDD 833 414 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=107760 $Y=59850 $D=111
M5754 426 476 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=114080 $Y=64310 $D=111
M5755 VDD 429 426 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=114560 $Y=64310 $D=111
M5756 838 448 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=114480 $Y=57110 $D=111
M5757 VDD 433 838 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=114960 $Y=57110 $D=111
M5758 430 443 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=116080 $Y=57110 $D=111
M5759 VDD 838 430 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=116560 $Y=57110 $D=111
M5760 439 443 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=117680 $Y=64310 $D=111
M5761 VDD 429 439 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=118160 $Y=64310 $D=111
M5762 427 477 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=121680 $Y=23850 $D=111
M5763 VDD 469 427 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=122160 $Y=23850 $D=111
M5764 477 456 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=122480 $Y=31050 $D=111
M5765 VDD 471 477 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=122960 $Y=31050 $D=111
M5766 844 457 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=123280 $Y=57110 $D=111
M5767 VDD 463 844 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=123760 $Y=57110 $D=111
M5768 481 844 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=126480 $Y=57110 $D=111
M5769 VDD 460 481 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=126960 $Y=57110 $D=111
M5770 520 502 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=132880 $Y=52650 $D=111
M5771 VDD 524 520 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=133360 $Y=52650 $D=111
M5772 519 515 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=133680 $Y=31050 $D=111
M5773 VDD 488 519 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=134160 $Y=31050 $D=111
M5774 560 559 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=138080 $Y=64310 $D=111
M5775 VDD 608 560 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=138560 $Y=64310 $D=111
M5776 522 558 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=140080 $Y=28310 $D=111
M5777 VDD 853 522 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=140560 $Y=28310 $D=111
M5778 854 548 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=143680 $Y=67050 $D=111
M5779 VDD 562 854 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=144160 $Y=67050 $D=111
M5780 557 601 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=147680 $Y=52650 $D=111
M5781 VDD 669 557 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=148160 $Y=52650 $D=111
M5782 626 602 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=149680 $Y=59850 $D=111
M5783 VDD 595 626 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=150160 $Y=59850 $D=111
M5784 614 609 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=154480 $Y=59850 $D=111
M5785 VDD 622 614 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=154960 $Y=59850 $D=111
M5786 624 625 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=157680 $Y=49910 $D=111
M5787 VDD 642 624 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=158160 $Y=49910 $D=111
M5788 633 632 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=161680 $Y=42710 $D=111
M5789 VDD 639 633 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=162160 $Y=42710 $D=111
M5790 692 617 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=164480 $Y=67050 $D=111
M5791 VDD 657 692 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=164960 $Y=67050 $D=111
M5792 712 710 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=166480 $Y=45450 $D=111
M5793 VDD 669 712 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=166960 $Y=45450 $D=111
M5794 679 576 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=166480 $Y=64310 $D=111
M5795 VDD 670 679 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=166960 $Y=64310 $D=111
M5796 676 724 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=166880 $Y=42710 $D=111
M5797 VDD 671 676 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=167360 $Y=42710 $D=111
M5798 713 685 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=167280 $Y=57110 $D=111
M5799 VDD 673 713 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=167760 $Y=57110 $D=111
M5800 724 726 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=167680 $Y=38250 $D=111
M5801 VDD 675 724 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=168160 $Y=38250 $D=111
M5802 695 684 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=170080 $Y=64310 $D=111
M5803 VDD 677 695 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=170560 $Y=64310 $D=111
M5804 785 696 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=171680 $Y=64310 $D=111
M5805 VDD 636 785 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=172160 $Y=64310 $D=111
M5806 863 732 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=173280 $Y=59850 $D=111
M5807 VDD 707 863 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=173760 $Y=59850 $D=111
M5808 735 683 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=174480 $Y=35510 $D=111
M5809 VDD 709 735 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=174960 $Y=35510 $D=111
M5810 715 723 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=175280 $Y=23850 $D=111
M5811 VDD 761 715 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=175760 $Y=23850 $D=111
M5812 736 652 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=175680 $Y=64310 $D=111
M5813 VDD 744 736 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=176160 $Y=64310 $D=111
M5814 723 717 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=176880 $Y=23850 $D=111
M5815 VDD 748 723 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=177360 $Y=23850 $D=111
M5816 752 749 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=179280 $Y=38250 $D=111
M5817 VDD 742 752 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=179760 $Y=38250 $D=111
M5818 865 759 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=182880 $Y=38250 $D=111
M5819 VDD 778 865 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=183360 $Y=38250 $D=111
M5820 VDD 10 1993 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=10810 $Y=13940 $D=111
M5821 1994 11 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=11440 $Y=13940 $D=111
M5822 798 1993 1994 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=11760 $Y=13940 $D=111
M5823 VDD 25 1995 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=12010 $Y=60160 $D=111
M5824 1996 23 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=12640 $Y=59620 $D=111
M5825 24 1995 1996 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=12960 $Y=59620 $D=111
M5826 VDD 41 1997 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=14010 $Y=60160 $D=111
M5827 1998 23 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=14640 $Y=59620 $D=111
M5828 18 1997 1998 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=14960 $Y=59620 $D=111
M5829 VDD 28 1999 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=14810 $Y=38560 $D=111
M5830 2000 23 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=15440 $Y=38020 $D=111
M5831 801 1999 2000 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=15760 $Y=38020 $D=111
M5832 VDD 122 2001 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=30010 $Y=16960 $D=111
M5833 2002 11 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=30640 $Y=16420 $D=111
M5834 95 2001 2002 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=30960 $Y=16420 $D=111
M5835 VDD 817 2003 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=59610 $Y=16960 $D=111
M5836 2004 11 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=60240 $Y=16420 $D=111
M5837 226 2003 2004 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=60560 $Y=16420 $D=111
M5838 VDD 257 2005 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=69610 $Y=21140 $D=111
M5839 2006 271 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=70240 $Y=21140 $D=111
M5840 261 2005 2006 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=70560 $Y=21140 $D=111
M5841 VDD 217 2007 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=71610 $Y=24160 $D=111
M5842 2008 148 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=72240 $Y=23620 $D=111
M5843 274 2007 2008 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=72560 $Y=23620 $D=111
M5844 VDD 826 2009 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=76810 $Y=21140 $D=111
M5845 2010 300 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=77440 $Y=21140 $D=111
M5846 827 2009 2010 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=77760 $Y=21140 $D=111
M5847 VDD 370 2011 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=104810 $Y=35540 $D=111
M5848 2012 409 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=105440 $Y=35540 $D=111
M5849 386 2011 2012 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=105760 $Y=35540 $D=111
M5850 VDD 573 2013 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=145610 $Y=31360 $D=111
M5851 2014 582 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=146240 $Y=30820 $D=111
M5852 577 2013 2014 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=146560 $Y=30820 $D=111
M5853 VDD 634 2015 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=153610 $Y=49940 $D=111
M5854 2016 592 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=154240 $Y=49940 $D=111
M5855 613 2015 2016 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=154560 $Y=49940 $D=111
M5856 VDD 663 2017 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=156010 $Y=42740 $D=111
M5857 2018 592 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=156640 $Y=42740 $D=111
M5858 647 2017 2018 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=156960 $Y=42740 $D=111
M5859 VDD 865 2019 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.01368e-13 as=9.6e-14 pd=7.10526e-07 ps=1.24e-06 nrd=1.12632 nrs=1.06667 sa=3.2e-07 sb=1.35e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=3.6e-15 panw8=0 panw9=0 panw10=0 $X=182810 $Y=28340 $D=111
M5860 2020 681 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.83832e-13 pd=1.04e-06 ps=1.98947e-06 nrd=0.119048 nrs=0.402256 sa=6.15714e-07 sb=7.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=183440 $Y=28340 $D=111
M5861 868 2019 2020 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.36e-13 as=8.4e-14 pd=2.48e-06 ps=1.04e-06 nrd=0.47619 nrs=0.119048 sa=9.35714e-07 sb=4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=183760 $Y=28340 $D=111
M5862 VDD 79 2022 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=25210 $Y=64310 $D=111
M5863 2022 79 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=25690 $Y=64310 $D=111
M5864 VDD 79 2022 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=26170 $Y=64310 $D=111
M5865 2021 110 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=26650 $Y=64310 $D=111
M5866 96 110 2022 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=27700 $Y=64530 $D=111
M5867 2022 110 96 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=28180 $Y=64530 $D=111
M5868 96 110 2022 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=28660 $Y=64530 $D=111
M5869 2023 2021 96 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=29140 $Y=64530 $D=111
M5870 96 2021 2023 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=29620 $Y=64530 $D=111
M5871 2023 2021 96 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=30100 $Y=64530 $D=111
M5872 VDD 2022 2023 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=30860 $Y=64310 $D=111
M5873 2023 2022 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=31340 $Y=64310 $D=111
M5874 VDD 2022 2023 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=31820 $Y=64310 $D=111
M5875 VDD 86 2025 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=25210 $Y=66650 $D=111
M5876 2025 86 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=25690 $Y=66650 $D=111
M5877 VDD 86 2025 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=26170 $Y=66650 $D=111
M5878 2024 79 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=26650 $Y=66470 $D=111
M5879 73 79 2025 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=27700 $Y=66430 $D=111
M5880 2025 79 73 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=28180 $Y=66430 $D=111
M5881 73 79 2025 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=28660 $Y=66430 $D=111
M5882 2026 2024 73 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=29140 $Y=66430 $D=111
M5883 73 2024 2026 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=29620 $Y=66430 $D=111
M5884 2026 2024 73 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=30100 $Y=66430 $D=111
M5885 VDD 2025 2026 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=30860 $Y=66650 $D=111
M5886 2026 2025 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=31340 $Y=66650 $D=111
M5887 VDD 2025 2026 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=31820 $Y=66650 $D=111
M5888 VDD 141 2028 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=38410 $Y=28310 $D=111
M5889 2028 141 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=38890 $Y=28310 $D=111
M5890 VDD 141 2028 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=39370 $Y=28310 $D=111
M5891 2027 163 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=39850 $Y=28310 $D=111
M5892 165 163 2028 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=40900 $Y=28530 $D=111
M5893 2028 163 165 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=41380 $Y=28530 $D=111
M5894 165 163 2028 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=41860 $Y=28530 $D=111
M5895 2029 2027 165 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=42340 $Y=28530 $D=111
M5896 165 2027 2029 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=42820 $Y=28530 $D=111
M5897 2029 2027 165 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=43300 $Y=28530 $D=111
M5898 VDD 2028 2029 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=44060 $Y=28310 $D=111
M5899 2029 2028 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=44540 $Y=28310 $D=111
M5900 VDD 2028 2029 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=45020 $Y=28310 $D=111
M5901 VDD 135 2031 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=39210 $Y=30650 $D=111
M5902 2031 135 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=39690 $Y=30650 $D=111
M5903 VDD 135 2031 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=40170 $Y=30650 $D=111
M5904 2030 123 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=40650 $Y=30470 $D=111
M5905 199 123 2031 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=41700 $Y=30430 $D=111
M5906 2031 123 199 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=42180 $Y=30430 $D=111
M5907 199 123 2031 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=42660 $Y=30430 $D=111
M5908 2032 2030 199 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=43140 $Y=30430 $D=111
M5909 199 2030 2032 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=43620 $Y=30430 $D=111
M5910 2032 2030 199 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=44100 $Y=30430 $D=111
M5911 VDD 2031 2032 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=44860 $Y=30650 $D=111
M5912 2032 2031 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=45340 $Y=30650 $D=111
M5913 VDD 2031 2032 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=45820 $Y=30650 $D=111
M5914 VDD 192 2034 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=44810 $Y=35510 $D=111
M5915 2034 192 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=45290 $Y=35510 $D=111
M5916 VDD 192 2034 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=45770 $Y=35510 $D=111
M5917 2033 163 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=46250 $Y=35510 $D=111
M5918 144 163 2034 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=47300 $Y=35730 $D=111
M5919 2034 163 144 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=47780 $Y=35730 $D=111
M5920 144 163 2034 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=48260 $Y=35730 $D=111
M5921 2035 2033 144 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=48740 $Y=35730 $D=111
M5922 144 2033 2035 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=49220 $Y=35730 $D=111
M5923 2035 2033 144 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=49700 $Y=35730 $D=111
M5924 VDD 2034 2035 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=50460 $Y=35510 $D=111
M5925 2035 2034 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=50940 $Y=35510 $D=111
M5926 VDD 2034 2035 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=51420 $Y=35510 $D=111
M5927 VDD 49 2037 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=47210 $Y=28310 $D=111
M5928 2037 49 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=47690 $Y=28310 $D=111
M5929 VDD 49 2037 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=48170 $Y=28310 $D=111
M5930 2036 113 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=48650 $Y=28310 $D=111
M5931 203 113 2037 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=49700 $Y=28530 $D=111
M5932 2037 113 203 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=50180 $Y=28530 $D=111
M5933 203 113 2037 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=50660 $Y=28530 $D=111
M5934 2038 2036 203 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=51140 $Y=28530 $D=111
M5935 203 2036 2038 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=51620 $Y=28530 $D=111
M5936 2038 2036 203 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=52100 $Y=28530 $D=111
M5937 VDD 2037 2038 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=52860 $Y=28310 $D=111
M5938 2038 2037 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=53340 $Y=28310 $D=111
M5939 VDD 2037 2038 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=53820 $Y=28310 $D=111
M5940 VDD 135 2040 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=55610 $Y=45050 $D=111
M5941 2040 135 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=56090 $Y=45050 $D=111
M5942 VDD 135 2040 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=56570 $Y=45050 $D=111
M5943 2039 123 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=57050 $Y=44870 $D=111
M5944 285 123 2040 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=58100 $Y=44830 $D=111
M5945 2040 123 285 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=58580 $Y=44830 $D=111
M5946 285 123 2040 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=59060 $Y=44830 $D=111
M5947 2041 2039 285 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=59540 $Y=44830 $D=111
M5948 285 2039 2041 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=60020 $Y=44830 $D=111
M5949 2041 2039 285 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=60500 $Y=44830 $D=111
M5950 VDD 2040 2041 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=61260 $Y=45050 $D=111
M5951 2041 2040 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=61740 $Y=45050 $D=111
M5952 VDD 2040 2041 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=62220 $Y=45050 $D=111
M5953 VDD 272 2043 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=60010 $Y=73850 $D=111
M5954 2043 272 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=60490 $Y=73850 $D=111
M5955 VDD 272 2043 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=60970 $Y=73850 $D=111
M5956 2042 268 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=61450 $Y=73670 $D=111
M5957 819 268 2043 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=62500 $Y=73630 $D=111
M5958 2043 268 819 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=62980 $Y=73630 $D=111
M5959 819 268 2043 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=63460 $Y=73630 $D=111
M5960 2044 2042 819 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=63940 $Y=73630 $D=111
M5961 819 2042 2044 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=64420 $Y=73630 $D=111
M5962 2044 2042 819 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=64900 $Y=73630 $D=111
M5963 VDD 2043 2044 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=65660 $Y=73850 $D=111
M5964 2044 2043 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=66140 $Y=73850 $D=111
M5965 VDD 2043 2044 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=66620 $Y=73850 $D=111
M5966 VDD 289 2046 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=60410 $Y=71510 $D=111
M5967 2046 289 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=60890 $Y=71510 $D=111
M5968 VDD 289 2046 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=61370 $Y=71510 $D=111
M5969 2045 819 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=61850 $Y=71510 $D=111
M5970 238 819 2046 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=62900 $Y=71730 $D=111
M5971 2046 819 238 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=63380 $Y=71730 $D=111
M5972 238 819 2046 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=63860 $Y=71730 $D=111
M5973 2047 2045 238 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=64340 $Y=71730 $D=111
M5974 238 2045 2047 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=64820 $Y=71730 $D=111
M5975 2047 2045 238 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=65300 $Y=71730 $D=111
M5976 VDD 2046 2047 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=66060 $Y=71510 $D=111
M5977 2047 2046 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=66540 $Y=71510 $D=111
M5978 VDD 2046 2047 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=67020 $Y=71510 $D=111
M5979 VDD 239 2049 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=65210 $Y=59450 $D=111
M5980 2049 239 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=65690 $Y=59450 $D=111
M5981 VDD 239 2049 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=66170 $Y=59450 $D=111
M5982 2048 248 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=66650 $Y=59270 $D=111
M5983 253 248 2049 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=67700 $Y=59230 $D=111
M5984 2049 248 253 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=68180 $Y=59230 $D=111
M5985 253 248 2049 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=68660 $Y=59230 $D=111
M5986 2050 2048 253 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=69140 $Y=59230 $D=111
M5987 253 2048 2050 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=69620 $Y=59230 $D=111
M5988 2050 2048 253 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=70100 $Y=59230 $D=111
M5989 VDD 2049 2050 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=70860 $Y=59450 $D=111
M5990 2050 2049 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=71340 $Y=59450 $D=111
M5991 VDD 2049 2050 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=71820 $Y=59450 $D=111
M5992 VDD 49 2052 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=67210 $Y=28310 $D=111
M5993 2052 49 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=67690 $Y=28310 $D=111
M5994 VDD 49 2052 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=68170 $Y=28310 $D=111
M5995 2051 170 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=68650 $Y=28310 $D=111
M5996 212 170 2052 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=69700 $Y=28530 $D=111
M5997 2052 170 212 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=70180 $Y=28530 $D=111
M5998 212 170 2052 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=70660 $Y=28530 $D=111
M5999 2053 2051 212 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=71140 $Y=28530 $D=111
M6000 212 2051 2053 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=71620 $Y=28530 $D=111
M6001 2053 2051 212 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=72100 $Y=28530 $D=111
M6002 VDD 2052 2053 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=72860 $Y=28310 $D=111
M6003 2053 2052 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=73340 $Y=28310 $D=111
M6004 VDD 2052 2053 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=73820 $Y=28310 $D=111
M6005 VDD 254 2055 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=67210 $Y=30650 $D=111
M6006 2055 254 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=67690 $Y=30650 $D=111
M6007 VDD 254 2055 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=68170 $Y=30650 $D=111
M6008 2054 170 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=68650 $Y=30470 $D=111
M6009 267 170 2055 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=69700 $Y=30430 $D=111
M6010 2055 170 267 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=70180 $Y=30430 $D=111
M6011 267 170 2055 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=70660 $Y=30430 $D=111
M6012 2056 2054 267 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=71140 $Y=30430 $D=111
M6013 267 2054 2056 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=71620 $Y=30430 $D=111
M6014 2056 2054 267 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=72100 $Y=30430 $D=111
M6015 VDD 2055 2056 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=72860 $Y=30650 $D=111
M6016 2056 2055 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=73340 $Y=30650 $D=111
M6017 VDD 2055 2056 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=73820 $Y=30650 $D=111
M6018 VDD 176 2058 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=79610 $Y=42710 $D=111
M6019 2058 176 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=80090 $Y=42710 $D=111
M6020 VDD 176 2058 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=80570 $Y=42710 $D=111
M6021 2057 307 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=81050 $Y=42710 $D=111
M6022 313 307 2058 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=82100 $Y=42930 $D=111
M6023 2058 307 313 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=82580 $Y=42930 $D=111
M6024 313 307 2058 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=83060 $Y=42930 $D=111
M6025 2059 2057 313 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=83540 $Y=42930 $D=111
M6026 313 2057 2059 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=84020 $Y=42930 $D=111
M6027 2059 2057 313 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=84500 $Y=42930 $D=111
M6028 VDD 2058 2059 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=85260 $Y=42710 $D=111
M6029 2059 2058 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=85740 $Y=42710 $D=111
M6030 VDD 2058 2059 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=86220 $Y=42710 $D=111
M6031 VDD 354 2061 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=98010 $Y=42710 $D=111
M6032 2061 354 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=98490 $Y=42710 $D=111
M6033 VDD 354 2061 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=98970 $Y=42710 $D=111
M6034 2060 367 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=99450 $Y=42710 $D=111
M6035 419 367 2061 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=100500 $Y=42930 $D=111
M6036 2061 367 419 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=100980 $Y=42930 $D=111
M6037 419 367 2061 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=101460 $Y=42930 $D=111
M6038 2062 2060 419 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=101940 $Y=42930 $D=111
M6039 419 2060 2062 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=102420 $Y=42930 $D=111
M6040 2062 2060 419 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=102900 $Y=42930 $D=111
M6041 VDD 2061 2062 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=103660 $Y=42710 $D=111
M6042 2062 2061 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=104140 $Y=42710 $D=111
M6043 VDD 2061 2062 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=104620 $Y=42710 $D=111
M6044 VDD 909 2064 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=98410 $Y=71510 $D=111
M6045 2064 909 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=98890 $Y=71510 $D=111
M6046 VDD 909 2064 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=99370 $Y=71510 $D=111
M6047 2063 383 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=99850 $Y=71510 $D=111
M6048 378 383 2064 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=100900 $Y=71730 $D=111
M6049 2064 383 378 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=101380 $Y=71730 $D=111
M6050 378 383 2064 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=101860 $Y=71730 $D=111
M6051 2065 2063 378 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=102340 $Y=71730 $D=111
M6052 378 2063 2065 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=102820 $Y=71730 $D=111
M6053 2065 2063 378 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=103300 $Y=71730 $D=111
M6054 VDD 2064 2065 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=104060 $Y=71510 $D=111
M6055 2065 2064 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=104540 $Y=71510 $D=111
M6056 VDD 2064 2065 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=105020 $Y=71510 $D=111
M6057 VDD 481 2067 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=121210 $Y=59450 $D=111
M6058 2067 481 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=121690 $Y=59450 $D=111
M6059 VDD 481 2067 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=122170 $Y=59450 $D=111
M6060 2066 464 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=122650 $Y=59270 $D=111
M6061 487 464 2067 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=123700 $Y=59230 $D=111
M6062 2067 464 487 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=124180 $Y=59230 $D=111
M6063 487 464 2067 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=124660 $Y=59230 $D=111
M6064 2068 2066 487 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=125140 $Y=59230 $D=111
M6065 487 2066 2068 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=125620 $Y=59230 $D=111
M6066 2068 2066 487 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=126100 $Y=59230 $D=111
M6067 VDD 2067 2068 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=126860 $Y=59450 $D=111
M6068 2068 2067 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=127340 $Y=59450 $D=111
M6069 VDD 2067 2068 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=127820 $Y=59450 $D=111
M6070 VDD 578 2070 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=144810 $Y=64310 $D=111
M6071 2070 578 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=145290 $Y=64310 $D=111
M6072 VDD 578 2070 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=145770 $Y=64310 $D=111
M6073 2069 583 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=146250 $Y=64310 $D=111
M6074 590 583 2070 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=147300 $Y=64530 $D=111
M6075 2070 583 590 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=147780 $Y=64530 $D=111
M6076 590 583 2070 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=148260 $Y=64530 $D=111
M6077 2071 2069 590 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=148740 $Y=64530 $D=111
M6078 590 2069 2071 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=149220 $Y=64530 $D=111
M6079 2071 2069 590 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=149700 $Y=64530 $D=111
M6080 VDD 2070 2071 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=150460 $Y=64310 $D=111
M6081 2071 2070 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=150940 $Y=64310 $D=111
M6082 VDD 2070 2071 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=151420 $Y=64310 $D=111
M6083 VDD 676 2073 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=168010 $Y=45050 $D=111
M6084 2073 676 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=168490 $Y=45050 $D=111
M6085 VDD 676 2073 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=168970 $Y=45050 $D=111
M6086 2072 702 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=169450 $Y=44870 $D=111
M6087 700 702 2073 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=170500 $Y=44830 $D=111
M6088 2073 702 700 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=170980 $Y=44830 $D=111
M6089 700 702 2073 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=171460 $Y=44830 $D=111
M6090 2074 2072 700 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=171940 $Y=44830 $D=111
M6091 700 2072 2074 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=172420 $Y=44830 $D=111
M6092 2074 2072 700 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=172900 $Y=44830 $D=111
M6093 VDD 2073 2074 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=173660 $Y=45050 $D=111
M6094 2074 2073 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=174140 $Y=45050 $D=111
M6095 VDD 2073 2074 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=174620 $Y=45050 $D=111
M6096 VDD 715 2076 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=181210 $Y=30650 $D=111
M6097 2076 715 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=181690 $Y=30650 $D=111
M6098 VDD 715 2076 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.95483e-13 as=1.872e-13 pd=1.45416e-06 ps=1.4e-06 nrd=0.180735 nrs=0.173077 sa=1.28e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=182170 $Y=30650 $D=111
M6099 2075 764 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.29317e-13 pd=3.08e-06 ps=1.70584e-06 nrd=0.262295 nrs=0.154069 sa=1.54164e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=182650 $Y=30470 $D=111
M6100 743 764 2076 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.328e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.307692 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=183700 $Y=30430 $D=111
M6101 2076 764 743 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=184180 $Y=30430 $D=111
M6102 743 764 2076 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.28e-06 sb=1.98942e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=184660 $Y=30430 $D=111
M6103 2077 2075 743 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.76e-06 sb=1.88788e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=185140 $Y=30430 $D=111
M6104 743 2075 2077 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=1.78635e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=185620 $Y=30430 $D=111
M6105 2077 2075 743 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.768e-13 as=1.872e-13 pd=1.9e-06 ps=1.4e-06 nrd=0.348373 nrs=0.173077 sa=2e-06 sb=1.68481e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=186100 $Y=30430 $D=111
M6106 VDD 2076 2077 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=3.768e-13 pd=1.4e-06 ps=1.9e-06 nrd=0.173077 nrs=0.348373 sa=1.68904e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=1.248e-13 $X=186860 $Y=30650 $D=111
M6107 2077 2076 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.79058e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.656e-13 panw10=0 $X=187340 $Y=30650 $D=111
M6108 VDD 2076 2077 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.307692 nrs=0.173077 sa=1.89212e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.488e-13 panw9=4.08e-14 panw10=0 $X=187820 $Y=30650 $D=111
M6109 2079 52 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=18940 $Y=30880 $D=111
M6110 VDD 52 2079 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=19420 $Y=30880 $D=111
M6111 2079 52 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=19900 $Y=30880 $D=111
M6112 VDD 52 2079 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=20380 $Y=30880 $D=111
M6113 2078 70 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=20920 $Y=30470 $D=111
M6114 26 70 2080 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=21740 $Y=30510 $D=111
M6115 2080 70 26 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=22220 $Y=30510 $D=111
M6116 26 70 2080 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=22700 $Y=30510 $D=111
M6117 2079 2078 26 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=23180 $Y=30510 $D=111
M6118 26 2078 2079 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=23660 $Y=30510 $D=111
M6119 2079 2078 26 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=24140 $Y=30510 $D=111
M6120 VDD 2079 2080 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=24960 $Y=30650 $D=111
M6121 2080 2079 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=25440 $Y=30650 $D=111
M6122 VDD 2079 2080 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=25920 $Y=30710 $D=111
M6123 2082 109 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=25340 $Y=52480 $D=111
M6124 VDD 109 2082 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=25820 $Y=52480 $D=111
M6125 2082 109 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=26300 $Y=52480 $D=111
M6126 VDD 109 2082 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=26780 $Y=52480 $D=111
M6127 2081 99 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=27320 $Y=52070 $D=111
M6128 92 99 2083 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=28140 $Y=52110 $D=111
M6129 2083 99 92 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=28620 $Y=52110 $D=111
M6130 92 99 2083 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=29100 $Y=52110 $D=111
M6131 2082 2081 92 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=29580 $Y=52110 $D=111
M6132 92 2081 2082 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=30060 $Y=52110 $D=111
M6133 2082 2081 92 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=30540 $Y=52110 $D=111
M6134 VDD 2082 2083 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=31360 $Y=52250 $D=111
M6135 2083 2082 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=31840 $Y=52250 $D=111
M6136 VDD 2082 2083 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=32320 $Y=52310 $D=111
M6137 2085 211 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=31740 $Y=57140 $D=111
M6138 VDD 211 2085 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=32220 $Y=57140 $D=111
M6139 2085 211 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=32700 $Y=57140 $D=111
M6140 VDD 211 2085 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=33180 $Y=57140 $D=111
M6141 2084 160 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=33720 $Y=57110 $D=111
M6142 99 160 2086 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=34540 $Y=57250 $D=111
M6143 2086 160 99 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=35020 $Y=57250 $D=111
M6144 99 160 2086 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=35500 $Y=57250 $D=111
M6145 2085 2084 99 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=35980 $Y=57250 $D=111
M6146 99 2084 2085 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=36460 $Y=57250 $D=111
M6147 2085 2084 99 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=36940 $Y=57250 $D=111
M6148 VDD 2085 2086 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=37760 $Y=57110 $D=111
M6149 2086 2085 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=38240 $Y=57110 $D=111
M6150 VDD 2085 2086 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=38720 $Y=57110 $D=111
M6151 2088 140 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=46540 $Y=21140 $D=111
M6152 VDD 140 2088 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=47020 $Y=21140 $D=111
M6153 2088 140 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=47500 $Y=21140 $D=111
M6154 VDD 140 2088 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=47980 $Y=21140 $D=111
M6155 2087 173 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=48520 $Y=21110 $D=111
M6156 188 173 2089 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=49340 $Y=21250 $D=111
M6157 2089 173 188 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=49820 $Y=21250 $D=111
M6158 188 173 2089 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=50300 $Y=21250 $D=111
M6159 2088 2087 188 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=50780 $Y=21250 $D=111
M6160 188 2087 2088 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=51260 $Y=21250 $D=111
M6161 2088 2087 188 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=51740 $Y=21250 $D=111
M6162 VDD 2088 2089 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=52560 $Y=21110 $D=111
M6163 2089 2088 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=53040 $Y=21110 $D=111
M6164 VDD 2088 2089 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=53520 $Y=21110 $D=111
M6165 2091 201 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=52940 $Y=49940 $D=111
M6166 VDD 201 2091 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=53420 $Y=49940 $D=111
M6167 2091 201 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=53900 $Y=49940 $D=111
M6168 VDD 201 2091 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=54380 $Y=49940 $D=111
M6169 2090 195 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=54920 $Y=49910 $D=111
M6170 213 195 2092 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=55740 $Y=50050 $D=111
M6171 2092 195 213 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=56220 $Y=50050 $D=111
M6172 213 195 2092 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=56700 $Y=50050 $D=111
M6173 2091 2090 213 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=57180 $Y=50050 $D=111
M6174 213 2090 2091 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=57660 $Y=50050 $D=111
M6175 2091 2090 213 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=58140 $Y=50050 $D=111
M6176 VDD 2091 2092 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=58960 $Y=49910 $D=111
M6177 2092 2091 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=59440 $Y=49910 $D=111
M6178 VDD 2091 2092 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=59920 $Y=49910 $D=111
M6179 2094 210 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=54140 $Y=59680 $D=111
M6180 VDD 210 2094 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=54620 $Y=59680 $D=111
M6181 2094 210 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=55100 $Y=59680 $D=111
M6182 VDD 210 2094 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=55580 $Y=59680 $D=111
M6183 2093 220 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=56120 $Y=59270 $D=111
M6184 230 220 2095 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=56940 $Y=59310 $D=111
M6185 2095 220 230 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=57420 $Y=59310 $D=111
M6186 230 220 2095 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=57900 $Y=59310 $D=111
M6187 2094 2093 230 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=58380 $Y=59310 $D=111
M6188 230 2093 2094 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=58860 $Y=59310 $D=111
M6189 2094 2093 230 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=59340 $Y=59310 $D=111
M6190 VDD 2094 2095 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=60160 $Y=59450 $D=111
M6191 2095 2094 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=60640 $Y=59450 $D=111
M6192 VDD 2094 2095 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=61120 $Y=59510 $D=111
M6193 2097 135 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=59340 $Y=28340 $D=111
M6194 VDD 135 2097 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=59820 $Y=28340 $D=111
M6195 2097 135 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=60300 $Y=28340 $D=111
M6196 VDD 135 2097 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=60780 $Y=28340 $D=111
M6197 2096 231 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=61320 $Y=28310 $D=111
M6198 236 231 2098 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=62140 $Y=28450 $D=111
M6199 2098 231 236 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=62620 $Y=28450 $D=111
M6200 236 231 2098 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=63100 $Y=28450 $D=111
M6201 2097 2096 236 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=63580 $Y=28450 $D=111
M6202 236 2096 2097 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=64060 $Y=28450 $D=111
M6203 2097 2096 236 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=64540 $Y=28450 $D=111
M6204 VDD 2097 2098 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=65360 $Y=28310 $D=111
M6205 2098 2097 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=65840 $Y=28310 $D=111
M6206 VDD 2097 2098 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=66320 $Y=28310 $D=111
M6207 2100 263 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=60140 $Y=38080 $D=111
M6208 VDD 263 2100 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=60620 $Y=38080 $D=111
M6209 2100 263 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=61100 $Y=38080 $D=111
M6210 VDD 263 2100 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=61580 $Y=38080 $D=111
M6211 2099 228 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=62120 $Y=37670 $D=111
M6212 237 228 2101 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=62940 $Y=37710 $D=111
M6213 2101 228 237 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=63420 $Y=37710 $D=111
M6214 237 228 2101 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=63900 $Y=37710 $D=111
M6215 2100 2099 237 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=64380 $Y=37710 $D=111
M6216 237 2099 2100 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=64860 $Y=37710 $D=111
M6217 2100 2099 237 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=65340 $Y=37710 $D=111
M6218 VDD 2100 2101 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=66160 $Y=37850 $D=111
M6219 2101 2100 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=66640 $Y=37850 $D=111
M6220 VDD 2100 2101 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=67120 $Y=37910 $D=111
M6221 2103 359 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=86940 $Y=57140 $D=111
M6222 VDD 359 2103 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=87420 $Y=57140 $D=111
M6223 2103 359 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=87900 $Y=57140 $D=111
M6224 VDD 359 2103 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=88380 $Y=57140 $D=111
M6225 2102 352 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=88920 $Y=57110 $D=111
M6226 355 352 2104 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=89740 $Y=57250 $D=111
M6227 2104 352 355 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=90220 $Y=57250 $D=111
M6228 355 352 2104 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=90700 $Y=57250 $D=111
M6229 2103 2102 355 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=91180 $Y=57250 $D=111
M6230 355 2102 2103 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=91660 $Y=57250 $D=111
M6231 2103 2102 355 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=92140 $Y=57250 $D=111
M6232 VDD 2103 2104 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=92960 $Y=57110 $D=111
M6233 2104 2103 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=93440 $Y=57110 $D=111
M6234 VDD 2103 2104 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=93920 $Y=57110 $D=111
M6235 2106 363 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=90940 $Y=52480 $D=111
M6236 VDD 363 2106 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=91420 $Y=52480 $D=111
M6237 2106 363 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=91900 $Y=52480 $D=111
M6238 VDD 363 2106 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=92380 $Y=52480 $D=111
M6239 2105 348 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=92920 $Y=52070 $D=111
M6240 352 348 2107 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=93740 $Y=52110 $D=111
M6241 2107 348 352 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=94220 $Y=52110 $D=111
M6242 352 348 2107 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=94700 $Y=52110 $D=111
M6243 2106 2105 352 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=95180 $Y=52110 $D=111
M6244 352 2105 2106 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=95660 $Y=52110 $D=111
M6245 2106 2105 352 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=96140 $Y=52110 $D=111
M6246 VDD 2106 2107 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=96960 $Y=52250 $D=111
M6247 2107 2106 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=97440 $Y=52250 $D=111
M6248 VDD 2106 2107 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=97920 $Y=52310 $D=111
M6249 2109 398 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=99340 $Y=52480 $D=111
M6250 VDD 398 2109 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=99820 $Y=52480 $D=111
M6251 2109 398 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=100300 $Y=52480 $D=111
M6252 VDD 398 2109 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=100780 $Y=52480 $D=111
M6253 2108 395 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=101320 $Y=52070 $D=111
M6254 380 395 2110 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=102140 $Y=52110 $D=111
M6255 2110 395 380 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=102620 $Y=52110 $D=111
M6256 380 395 2110 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=103100 $Y=52110 $D=111
M6257 2109 2108 380 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=103580 $Y=52110 $D=111
M6258 380 2108 2109 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=104060 $Y=52110 $D=111
M6259 2109 2108 380 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=104540 $Y=52110 $D=111
M6260 VDD 2109 2110 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=105360 $Y=52250 $D=111
M6261 2110 2109 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=105840 $Y=52250 $D=111
M6262 VDD 2109 2110 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=106320 $Y=52310 $D=111
M6263 2112 426 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=108940 $Y=59680 $D=111
M6264 VDD 426 2112 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=109420 $Y=59680 $D=111
M6265 2112 426 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=109900 $Y=59680 $D=111
M6266 VDD 426 2112 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=110380 $Y=59680 $D=111
M6267 2111 415 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=110920 $Y=59270 $D=111
M6268 394 415 2113 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=111740 $Y=59310 $D=111
M6269 2113 415 394 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=112220 $Y=59310 $D=111
M6270 394 415 2113 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=112700 $Y=59310 $D=111
M6271 2112 2111 394 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=113180 $Y=59310 $D=111
M6272 394 2111 2112 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=113660 $Y=59310 $D=111
M6273 2112 2111 394 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=114140 $Y=59310 $D=111
M6274 VDD 2112 2113 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=114960 $Y=59450 $D=111
M6275 2113 2112 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=115440 $Y=59450 $D=111
M6276 VDD 2112 2113 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=115920 $Y=59510 $D=111
M6277 2115 507 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=125340 $Y=23680 $D=111
M6278 VDD 507 2115 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=125820 $Y=23680 $D=111
M6279 2115 507 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=126300 $Y=23680 $D=111
M6280 VDD 507 2115 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=126780 $Y=23680 $D=111
M6281 2114 483 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=127320 $Y=23270 $D=111
M6282 514 483 2116 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=128140 $Y=23310 $D=111
M6283 2116 483 514 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=128620 $Y=23310 $D=111
M6284 514 483 2116 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=129100 $Y=23310 $D=111
M6285 2115 2114 514 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=129580 $Y=23310 $D=111
M6286 514 2114 2115 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=130060 $Y=23310 $D=111
M6287 2115 2114 514 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=130540 $Y=23310 $D=111
M6288 VDD 2115 2116 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=131360 $Y=23450 $D=111
M6289 2116 2115 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=131840 $Y=23450 $D=111
M6290 VDD 2115 2116 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=132320 $Y=23510 $D=111
M6291 2118 498 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=128940 $Y=59680 $D=111
M6292 VDD 498 2118 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=129420 $Y=59680 $D=111
M6293 2118 498 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=129900 $Y=59680 $D=111
M6294 VDD 498 2118 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=130380 $Y=59680 $D=111
M6295 2117 511 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=130920 $Y=59270 $D=111
M6296 521 511 2119 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=131740 $Y=59310 $D=111
M6297 2119 511 521 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=132220 $Y=59310 $D=111
M6298 521 511 2119 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=132700 $Y=59310 $D=111
M6299 2118 2117 521 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=133180 $Y=59310 $D=111
M6300 521 2117 2118 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=133660 $Y=59310 $D=111
M6301 2118 2117 521 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=134140 $Y=59310 $D=111
M6302 VDD 2118 2119 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=134960 $Y=59450 $D=111
M6303 2119 2118 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=135440 $Y=59450 $D=111
M6304 VDD 2118 2119 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=135920 $Y=59510 $D=111
M6305 2121 555 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=137340 $Y=35540 $D=111
M6306 VDD 555 2121 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=137820 $Y=35540 $D=111
M6307 2121 555 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=138300 $Y=35540 $D=111
M6308 VDD 555 2121 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=138780 $Y=35540 $D=111
M6309 2120 542 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=139320 $Y=35510 $D=111
M6310 535 542 2122 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=140140 $Y=35650 $D=111
M6311 2122 542 535 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=140620 $Y=35650 $D=111
M6312 535 542 2122 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=141100 $Y=35650 $D=111
M6313 2121 2120 535 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=141580 $Y=35650 $D=111
M6314 535 2120 2121 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=142060 $Y=35650 $D=111
M6315 2121 2120 535 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=142540 $Y=35650 $D=111
M6316 VDD 2121 2122 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=143360 $Y=35510 $D=111
M6317 2122 2121 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=143840 $Y=35510 $D=111
M6318 VDD 2121 2122 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=144320 $Y=35510 $D=111
M6319 2124 672 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=156140 $Y=71540 $D=111
M6320 VDD 672 2124 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=156620 $Y=71540 $D=111
M6321 2124 672 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=157100 $Y=71540 $D=111
M6322 VDD 672 2124 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=157580 $Y=71540 $D=111
M6323 2123 857 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=158120 $Y=71510 $D=111
M6324 644 857 2125 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=158940 $Y=71650 $D=111
M6325 2125 857 644 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=159420 $Y=71650 $D=111
M6326 644 857 2125 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=159900 $Y=71650 $D=111
M6327 2124 2123 644 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=160380 $Y=71650 $D=111
M6328 644 2123 2124 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=160860 $Y=71650 $D=111
M6329 2124 2123 644 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=161340 $Y=71650 $D=111
M6330 VDD 2124 2125 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=162160 $Y=71510 $D=111
M6331 2125 2124 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=162640 $Y=71510 $D=111
M6332 VDD 2124 2125 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=163120 $Y=71510 $D=111
M6333 2127 861 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=169340 $Y=74080 $D=111
M6334 VDD 861 2127 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=169820 $Y=74080 $D=111
M6335 2127 861 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=170300 $Y=74080 $D=111
M6336 VDD 861 2127 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=170780 $Y=74080 $D=111
M6337 2126 763 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=171320 $Y=73670 $D=111
M6338 705 763 2128 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=172140 $Y=73710 $D=111
M6339 2128 763 705 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=172620 $Y=73710 $D=111
M6340 705 763 2128 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=173100 $Y=73710 $D=111
M6341 2127 2126 705 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=173580 $Y=73710 $D=111
M6342 705 2126 2127 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=174060 $Y=73710 $D=111
M6343 2127 2126 705 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=174540 $Y=73710 $D=111
M6344 VDD 2127 2128 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=175360 $Y=73850 $D=111
M6345 2128 2127 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=175840 $Y=73850 $D=111
M6346 VDD 2127 2128 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=176320 $Y=73910 $D=111
M6347 2130 774 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=179740 $Y=21140 $D=111
M6348 VDD 774 2130 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=180220 $Y=21140 $D=111
M6349 2130 774 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=180700 $Y=21140 $D=111
M6350 VDD 774 2130 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=181180 $Y=21140 $D=111
M6351 2129 787 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=181720 $Y=21110 $D=111
M6352 767 787 2131 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=182540 $Y=21250 $D=111
M6353 2131 787 767 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=183020 $Y=21250 $D=111
M6354 767 787 2131 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=183500 $Y=21250 $D=111
M6355 2130 2129 767 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=183980 $Y=21250 $D=111
M6356 767 2129 2130 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=184460 $Y=21250 $D=111
M6357 2130 2129 767 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=184940 $Y=21250 $D=111
M6358 VDD 2130 2131 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=185760 $Y=21110 $D=111
M6359 2131 2130 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=186240 $Y=21110 $D=111
M6360 VDD 2130 2131 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=9.8e-14 $X=186720 $Y=21110 $D=111
M6361 2133 753 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=180940 $Y=57140 $D=111
M6362 VDD 753 2133 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=181420 $Y=57140 $D=111
M6363 2133 753 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=181900 $Y=57140 $D=111
M6364 VDD 753 2133 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=182380 $Y=57140 $D=111
M6365 2132 866 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=182920 $Y=57110 $D=111
M6366 768 866 2134 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=183740 $Y=57250 $D=111
M6367 2134 866 768 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=184220 $Y=57250 $D=111
M6368 768 866 2134 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=184700 $Y=57250 $D=111
M6369 2133 2132 768 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=185180 $Y=57250 $D=111
M6370 768 2132 2133 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=185660 $Y=57250 $D=111
M6371 2133 2132 768 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=186140 $Y=57250 $D=111
M6372 VDD 2133 2134 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=1.248e-13 $X=186960 $Y=57110 $D=111
M6373 2134 2133 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.656e-13 panw10=0 $X=187440 $Y=57110 $D=111
M6374 VDD 2133 2134 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.22e-13 panw8=4.36e-14 panw9=3.36e-14 panw10=0 $X=187920 $Y=57110 $D=111
M6375 2136 738 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=3.63215e-13 pd=1.14e-06 ps=2.79623e-06 nrd=0.230769 nrs=0.597 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=180940 $Y=64340 $D=111
M6376 VDD 738 2136 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=8.4e-07 sb=1.73846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=181420 $Y=64340 $D=111
M6377 2136 738 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.404e-13 pd=1.14e-06 ps=1.14e-06 nrd=0.230769 nrs=0.230769 sa=1.32e-06 sb=1.25846e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=181900 $Y=64340 $D=111
M6378 VDD 738 2136 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85968e-13 as=1.404e-13 pd=1.30684e-06 ps=1.14e-06 nrd=0.305668 nrs=0.230769 sa=1.8e-06 sb=7.78462e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.32e-14 panw10=0 $X=182380 $Y=64340 $D=111
M6379 2135 751 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.776e-13 as=2.90874e-13 pd=3.08e-06 ps=2.04404e-06 nrd=0.186509 nrs=0.195427 sa=1.39836e-06 sb=2.27541e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.44e-14 $X=182920 $Y=64310 $D=111
M6380 777 751 2137 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=183740 $Y=64450 $D=111
M6381 2137 751 777 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=7.12308e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=184220 $Y=64450 $D=111
M6382 777 751 2137 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.19231e-06 sb=1.72308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=184700 $Y=64450 $D=111
M6383 2136 2135 777 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=1.67231e-06 sb=1.24308e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=185180 $Y=64450 $D=111
M6384 777 2135 2136 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.872e-13 pd=1.4e-06 ps=1.4e-06 nrd=0.173077 nrs=0.173077 sa=2e-06 sb=7.63077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=185660 $Y=64450 $D=111
M6385 2136 2135 777 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=1.872e-13 pd=2.72e-06 ps=1.4e-06 nrd=0.272189 nrs=0.173077 sa=2e-06 sb=2.83077e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=186140 $Y=64450 $D=111
M6386 VDD 2136 2137 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=2.416e-13 pd=1.4e-06 ps=2.72e-06 nrd=0.173077 nrs=0.223373 sa=2.32308e-07 sb=1.17e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=1.248e-13 $X=186960 $Y=64310 $D=111
M6387 2137 2136 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.87818e-13 as=1.872e-13 pd=1.44158e-06 ps=1.4e-06 nrd=0.173648 nrs=0.173077 sa=7.12308e-07 sb=6.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.656e-13 panw10=0 $X=187440 $Y=64310 $D=111
M6388 VDD 2136 2137 VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.82489e-13 as=1.76982e-13 pd=3.00222e-06 ps=1.35842e-06 nrd=0.294137 nrs=0.18428 sa=1.19429e-06 sb=2.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.22e-13 panw8=4.36e-14 panw9=3.36e-14 panw10=0 $X=187920 $Y=64310 $D=111
M6389 33 27 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=14550 $Y=28350 $D=111
M6390 VDD 62 33 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=15030 $Y=28350 $D=111
M6391 40 39 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=16150 $Y=21150 $D=111
M6392 VDD 133 40 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=16630 $Y=21150 $D=111
M6393 105 803 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=21750 $Y=71550 $D=111
M6394 VDD 65 105 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=22230 $Y=71550 $D=111
M6395 85 69 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=23750 $Y=66390 $D=111
M6396 VDD 121 85 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=24230 $Y=66390 $D=111
M6397 108 145 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=26550 $Y=37590 $D=111
M6398 VDD 87 108 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=27030 $Y=37590 $D=111
M6399 807 109 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=32950 $Y=59190 $D=111
M6400 VDD 138 807 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=33430 $Y=59190 $D=111
M6401 890 139 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=33750 $Y=66390 $D=111
M6402 VDD 138 890 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=34230 $Y=66390 $D=111
M6403 91 238 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=35350 $Y=71550 $D=111
M6404 VDD 191 91 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=35830 $Y=71550 $D=111
M6405 132 130 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=36550 $Y=21150 $D=111
M6406 VDD 125 132 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=37030 $Y=21150 $D=111
M6407 161 139 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=39750 $Y=64350 $D=111
M6408 VDD 109 161 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=40230 $Y=64350 $D=111
M6409 815 167 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=56550 $Y=21150 $D=111
M6410 VDD 205 815 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=57030 $Y=21150 $D=111
M6411 233 230 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=62550 $Y=59190 $D=111
M6412 VDD 818 233 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=63030 $Y=59190 $D=111
M6413 904 823 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=68950 $Y=71550 $D=111
M6414 VDD 821 904 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=69430 $Y=71550 $D=111
M6415 361 323 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=90950 $Y=73590 $D=111
M6416 VDD 342 361 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=91430 $Y=73590 $D=111
M6417 375 363 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=98950 $Y=57150 $D=111
M6418 VDD 360 375 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=99430 $Y=57150 $D=111
M6419 379 359 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=101350 $Y=59190 $D=111
M6420 VDD 360 379 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=101830 $Y=59190 $D=111
M6421 432 433 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=116150 $Y=64350 $D=111
M6422 VDD 448 432 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=116630 $Y=64350 $D=111
M6423 445 441 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=118150 $Y=30390 $D=111
M6424 VDD 450 445 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=118630 $Y=30390 $D=111
M6425 502 480 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=127750 $Y=42750 $D=111
M6426 VDD 845 502 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=128230 $Y=42750 $D=111
M6427 517 470 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=129750 $Y=42750 $D=111
M6428 VDD 493 517 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=130230 $Y=42750 $D=111
M6429 512 525 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=137750 $Y=44790 $D=111
M6430 VDD 510 512 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=138230 $Y=44790 $D=111
M6431 585 571 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=145750 $Y=35550 $D=111
M6432 VDD 577 585 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=146230 $Y=35550 $D=111
M6433 580 587 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=148550 $Y=49950 $D=111
M6434 VDD 613 580 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=149030 $Y=49950 $D=111
M6435 649 637 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=161750 $Y=49950 $D=111
M6436 VDD 647 649 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=162230 $Y=49950 $D=111
M6437 779 752 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.268e-13 as=4.32982e-13 pd=1.62e-06 ps=3.09273e-06 nrd=0.142857 nrs=0.272727 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=181350 $Y=37590 $D=111
M6438 VDD 781 779 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.268e-13 pd=3.09273e-06 ps=1.62e-06 nrd=0.272727 nrs=0.142857 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=181830 $Y=37590 $D=111
M6439 51 80 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=20920 $Y=64310 $D=111
M6440 54 51 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=19280 $Y=64310 $D=111
M6441 VDD 50 54 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=19760 $Y=64310 $D=111
M6442 847 504 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=129720 $Y=28310 $D=111
M6443 504 474 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=128080 $Y=28310 $D=111
M6444 VDD 486 504 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=128560 $Y=28310 $D=111
M6445 851 527 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=134520 $Y=28310 $D=111
M6446 509 501 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=132880 $Y=28310 $D=111
M6447 VDD 469 509 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=133360 $Y=28310 $D=111
M6448 853 528 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=138920 $Y=28310 $D=111
M6449 536 505 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=137280 $Y=28310 $D=111
M6450 VDD 529 536 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=137760 $Y=28310 $D=111
M6451 569 632 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=146520 $Y=28310 $D=111
M6452 554 568 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=144880 $Y=28310 $D=111
M6453 VDD 569 554 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=145360 $Y=28310 $D=111
M6454 595 581 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=148520 $Y=59850 $D=111
M6455 578 607 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=146880 $Y=59850 $D=111
M6456 VDD 595 578 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=147360 $Y=59850 $D=111
M6457 588 609 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=151720 $Y=57110 $D=111
M6458 607 597 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=150080 $Y=57110 $D=111
M6459 VDD 588 607 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=150560 $Y=57110 $D=111
M6460 629 660 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=163320 $Y=45450 $D=111
M6461 660 646 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=161680 $Y=45450 $D=111
M6462 VDD 630 660 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=162160 $Y=45450 $D=111
M6463 744 746 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.24e-13 pd=1.92e-06 ps=1.98e-06 nrd=0.5 nrs=0.546875 sa=3.5e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=181720 $Y=52650 $D=111
M6464 734 746 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=3.41426e-13 pd=1e-06 ps=2.68522e-06 nrd=0.28125 nrs=0.83356 sa=3.6e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=180080 $Y=52650 $D=111
M6465 VDD 750 734 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=1.152e-13 pd=2e-06 ps=1e-06 nrd=0.5625 nrs=0.28125 sa=8.4e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=180560 $Y=52650 $D=111
M6466 2197 26 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.092e-13 as=3.15467e-13 pd=9.5e-07 ps=2.52e-06 nrd=0.348214 nrs=1.00595 sa=3.6e-07 sb=1.99e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=11130 $Y=28350 $D=111
M6467 VDD 47 2197 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.56053e-13 as=1.092e-13 pd=1.06133e-06 ps=9.5e-07 nrd=0.497619 nrs=0.348214 sa=8.7e-07 sb=1.48e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=11640 $Y=28350 $D=111
M6468 66 2197 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.646e-13 as=3.5112e-13 pd=1.68e-06 ps=2.388e-06 nrd=0.166667 nrs=0.221164 sa=8.44444e-07 sb=9e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=12220 $Y=28350 $D=111
M6469 VDD 33 66 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.646e-13 pd=3.09273e-06 ps=1.68e-06 nrd=0.272727 nrs=0.166667 sa=1.38444e-06 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=12760 $Y=28350 $D=111
M6470 2201 151 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.092e-13 as=3.15467e-13 pd=9.5e-07 ps=2.52e-06 nrd=0.348214 nrs=1.00595 sa=3.6e-07 sb=1.99e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=51130 $Y=59890 $D=111
M6471 VDD 189 2201 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.56053e-13 as=1.092e-13 pd=1.06133e-06 ps=9.5e-07 nrd=0.497619 nrs=0.348214 sa=8.7e-07 sb=1.48e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=51640 $Y=59890 $D=111
M6472 340 2201 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.646e-13 as=3.5112e-13 pd=1.68e-06 ps=2.388e-06 nrd=0.166667 nrs=0.221164 sa=8.44444e-07 sb=9e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=52220 $Y=59190 $D=111
M6473 VDD 193 340 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.646e-13 pd=3.09273e-06 ps=1.68e-06 nrd=0.272727 nrs=0.166667 sa=1.38444e-06 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=52760 $Y=59190 $D=111
M6474 2205 215 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.092e-13 as=3.15467e-13 pd=9.5e-07 ps=2.52e-06 nrd=0.348214 nrs=1.00595 sa=3.6e-07 sb=1.99e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=62730 $Y=57150 $D=111
M6475 VDD 220 2205 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.56053e-13 as=1.092e-13 pd=1.06133e-06 ps=9.5e-07 nrd=0.497619 nrs=0.348214 sa=8.7e-07 sb=1.48e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=63240 $Y=57150 $D=111
M6476 275 2205 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.646e-13 as=3.5112e-13 pd=1.68e-06 ps=2.388e-06 nrd=0.166667 nrs=0.221164 sa=8.44444e-07 sb=9e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=63820 $Y=57150 $D=111
M6477 VDD 229 275 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.646e-13 pd=3.09273e-06 ps=1.68e-06 nrd=0.272727 nrs=0.166667 sa=1.38444e-06 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=64360 $Y=57150 $D=111
M6478 2209 268 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.092e-13 as=3.15467e-13 pd=9.5e-07 ps=2.52e-06 nrd=0.348214 nrs=1.00595 sa=3.6e-07 sb=1.99e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=71930 $Y=74290 $D=111
M6479 VDD 272 2209 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.56053e-13 as=1.092e-13 pd=1.06133e-06 ps=9.5e-07 nrd=0.497619 nrs=0.348214 sa=8.7e-07 sb=1.48e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=72440 $Y=74290 $D=111
M6480 308 2209 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.646e-13 as=3.5112e-13 pd=1.68e-06 ps=2.388e-06 nrd=0.166667 nrs=0.221164 sa=8.44444e-07 sb=9e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=73020 $Y=73590 $D=111
M6481 VDD 277 308 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.646e-13 pd=3.09273e-06 ps=1.68e-06 nrd=0.272727 nrs=0.166667 sa=1.38444e-06 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=73560 $Y=73590 $D=111
M6482 2213 761 VDD VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.092e-13 as=3.15467e-13 pd=9.5e-07 ps=2.52e-06 nrd=0.348214 nrs=1.00595 sa=3.6e-07 sb=1.99e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=179930 $Y=28350 $D=111
M6483 VDD 741 2213 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.56053e-13 as=1.092e-13 pd=1.06133e-06 ps=9.5e-07 nrd=0.497619 nrs=0.348214 sa=8.7e-07 sb=1.48e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-14 panw9=0 panw10=0 $X=180440 $Y=28350 $D=111
M6484 780 2213 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.646e-13 as=3.5112e-13 pd=1.68e-06 ps=2.388e-06 nrd=0.166667 nrs=0.221164 sa=8.44444e-07 sb=9e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=181020 $Y=28350 $D=111
M6485 VDD 756 780 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.32982e-13 as=2.646e-13 pd=3.09273e-06 ps=1.68e-06 nrd=0.272727 nrs=0.166667 sa=1.38444e-06 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=181560 $Y=28350 $D=111
M6486 2217 853 VDD VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=1.7e-13 pd=1.53e-06 ps=1.68e-06 nrd=0.576 nrs=0.68 sa=3.4e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=141670 $Y=28310 $D=111
M6487 VDD 536 2217 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.27697e-13 as=1.44e-13 pd=9.49438e-07 ps=1.53e-06 nrd=0.510787 nrs=0.576 sa=7.8e-07 sb=8.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=142110 $Y=28310 $D=111
M6488 555 2217 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=3.26903e-13 pd=3.2e-06 ps=2.43056e-06 nrd=0.25 nrs=0.199526 sa=7.06719e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=142640 $Y=28310 $D=111
M6489 2219 602 VDD VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=1.7e-13 pd=1.53e-06 ps=1.68e-06 nrd=0.576 nrs=0.68 sa=3.4e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=152470 $Y=64310 $D=111
M6490 VDD 614 2219 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.27697e-13 as=1.44e-13 pd=9.49438e-07 ps=1.53e-06 nrd=0.510787 nrs=0.576 sa=7.8e-07 sb=8.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=152910 $Y=64310 $D=111
M6491 608 2219 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=3.26903e-13 pd=3.2e-06 ps=2.43056e-06 nrd=0.25 nrs=0.199526 sa=7.06719e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=153440 $Y=64310 $D=111
M6492 2221 720 VDD VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=1.7e-13 pd=1.53e-06 ps=1.68e-06 nrd=0.576 nrs=0.68 sa=3.4e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=177270 $Y=38390 $D=111
M6493 VDD 735 2221 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.27697e-13 as=1.44e-13 pd=9.49438e-07 ps=1.53e-06 nrd=0.510787 nrs=0.576 sa=7.8e-07 sb=8.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=177710 $Y=38390 $D=111
M6494 778 2221 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=3.26903e-13 pd=3.2e-06 ps=2.43056e-06 nrd=0.25 nrs=0.199526 sa=7.06719e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=178240 $Y=37610 $D=111
M6495 2223 732 VDD VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=1.7e-13 pd=1.53e-06 ps=1.68e-06 nrd=0.576 nrs=0.68 sa=3.4e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=177670 $Y=57110 $D=111
M6496 VDD 734 2223 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.27697e-13 as=1.44e-13 pd=9.49438e-07 ps=1.53e-06 nrd=0.510787 nrs=0.576 sa=7.8e-07 sb=8.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=178110 $Y=57110 $D=111
M6497 753 2223 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=3.26903e-13 pd=3.2e-06 ps=2.43056e-06 nrd=0.25 nrs=0.199526 sa=7.06719e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=178640 $Y=57110 $D=111
M6498 2225 737 VDD VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=1.7e-13 pd=1.53e-06 ps=1.68e-06 nrd=0.576 nrs=0.68 sa=3.4e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=178470 $Y=23990 $D=111
M6499 VDD 761 2225 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.27697e-13 as=1.44e-13 pd=9.49438e-07 ps=1.53e-06 nrd=0.510787 nrs=0.576 sa=7.8e-07 sb=8.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=178910 $Y=23990 $D=111
M6500 755 2225 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=3.26903e-13 pd=3.2e-06 ps=2.43056e-06 nrd=0.25 nrs=0.199526 sa=7.06719e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=179440 $Y=23210 $D=111
M6501 2228 666 VDD VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.28e-14 as=3.334e-13 pd=6.8e-07 ps=2.9e-06 nrd=0.272727 nrs=1.72211 sa=3.5e-07 sb=1.21455e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=162840 $Y=52790 $D=111
M6502 650 659 2228 VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.92279e-14 as=5.28e-14 pd=8.59535e-07 ps=6.8e-07 nrd=0.460888 nrs=0.272727 sa=7.1e-07 sb=8.54545e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=163200 $Y=52790 $D=111
M6503 VDD 633 650 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.492e-13 as=8.51721e-14 pd=2.26e-06 ps=8.20465e-07 nrd=1.4127 nrs=0.482835 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=163720 $Y=52810 $D=111
M6504 2230 863 VDD VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.28e-14 as=3.334e-13 pd=6.8e-07 ps=2.9e-06 nrd=0.272727 nrs=1.72211 sa=3.5e-07 sb=1.21455e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=174440 $Y=57170 $D=111
M6505 718 725 2230 VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.92279e-14 as=5.28e-14 pd=8.59535e-07 ps=6.8e-07 nrd=0.460888 nrs=0.272727 sa=7.1e-07 sb=8.54545e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=174800 $Y=57170 $D=111
M6506 VDD 714 718 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.492e-13 as=8.51721e-14 pd=2.26e-06 ps=8.20465e-07 nrd=1.4127 nrs=0.482835 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=175320 $Y=57170 $D=111
M6507 2232 713 VDD VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.28e-14 as=3.334e-13 pd=6.8e-07 ps=2.9e-06 nrd=0.272727 nrs=1.72211 sa=3.5e-07 sb=1.21455e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=178040 $Y=52790 $D=111
M6508 739 659 2232 VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.92279e-14 as=5.28e-14 pd=8.59535e-07 ps=6.8e-07 nrd=0.460888 nrs=0.272727 sa=7.1e-07 sb=8.54545e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=178400 $Y=52790 $D=111
M6509 VDD 721 739 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.492e-13 as=8.51721e-14 pd=2.26e-06 ps=8.20465e-07 nrd=1.4127 nrs=0.482835 sa=1.23e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=178920 $Y=52810 $D=111
M6510 VDD clk 2233 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=4.08e-14 panw10=0 $X=9330 $Y=64310 $D=111
M6511 2241 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=1.176e-13 $X=9730 $Y=64310 $D=111
M6512 2235 2238 2241 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=10130 $Y=64310 $D=111
M6513 VDD 2233 2238 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=11070 $Y=64450 $D=111
M6514 2234 18 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=11470 $Y=64450 $D=111
M6515 2242 2238 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=12390 $Y=64590 $D=111
M6516 2236 2234 2242 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=12710 $Y=64590 $D=111
M6517 2244 2235 2236 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=13240 $Y=64490 $D=111
M6518 VDD 2237 2244 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=13560 $Y=64490 $D=111
M6519 2237 2236 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=13960 $Y=64490 $D=111
M6520 VDD 2236 2237 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=14440 $Y=64490 $D=111
M6521 2237 32 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=14880 $Y=64490 $D=111
M6522 2240 2235 2237 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=15360 $Y=64490 $D=111
M6523 2237 2235 2240 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=15840 $Y=64490 $D=111
M6524 2249 2239 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=16700 $Y=65010 $D=111
M6525 2240 2238 2249 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=17020 $Y=65010 $D=111
M6526 VDD 32 2240 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=17500 $Y=65010 $D=111
M6527 VDD 2240 2239 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=17820 $Y=64310 $D=111
M6528 260 2240 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=18220 $Y=64310 $D=111
M6529 VDD clk 2250 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=96530 $Y=31350 $D=111
M6530 2258 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=96930 $Y=30710 $D=111
M6531 2252 2255 2258 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=97330 $Y=30950 $D=111
M6532 VDD 2250 2255 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=98270 $Y=30390 $D=111
M6533 2251 386 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=98670 $Y=31190 $D=111
M6534 2259 2255 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=99590 $Y=30390 $D=111
M6535 2253 2251 2259 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=99910 $Y=30390 $D=111
M6536 2261 2252 2253 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=100440 $Y=31230 $D=111
M6537 VDD 2254 2261 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=100760 $Y=31230 $D=111
M6538 2254 2253 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=101160 $Y=30710 $D=111
M6539 VDD 2253 2254 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=101640 $Y=30710 $D=111
M6540 2254 374 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=102080 $Y=31110 $D=111
M6541 2257 2252 2254 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=102560 $Y=30770 $D=111
M6542 2254 2252 2257 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=103040 $Y=30710 $D=111
M6543 2266 2256 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=103900 $Y=30710 $D=111
M6544 2257 2255 2266 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=104220 $Y=30710 $D=111
M6545 VDD 374 2257 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=104700 $Y=30590 $D=111
M6546 VDD 2257 2256 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=105020 $Y=31410 $D=111
M6547 363 2257 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=105420 $Y=30390 $D=111
M6548 VDD clk 2267 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=109330 $Y=21110 $D=111
M6549 2275 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=109730 $Y=21110 $D=111
M6550 2269 2272 2275 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=110130 $Y=21110 $D=111
M6551 VDD 2267 2272 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=111070 $Y=21250 $D=111
M6552 2268 834 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=111470 $Y=21250 $D=111
M6553 2276 2272 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=112390 $Y=21390 $D=111
M6554 2270 2268 2276 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=112710 $Y=21390 $D=111
M6555 2278 2269 2270 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=113240 $Y=21290 $D=111
M6556 VDD 2271 2278 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=113560 $Y=21290 $D=111
M6557 2271 2270 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=113960 $Y=21290 $D=111
M6558 VDD 2270 2271 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=114440 $Y=21290 $D=111
M6559 2271 425 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=114880 $Y=21290 $D=111
M6560 2274 2269 2271 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=115360 $Y=21290 $D=111
M6561 2271 2269 2274 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=115840 $Y=21290 $D=111
M6562 2283 2273 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=116700 $Y=21810 $D=111
M6563 2274 2272 2283 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=117020 $Y=21810 $D=111
M6564 VDD 425 2274 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=117500 $Y=21810 $D=111
M6565 VDD 2274 2273 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=117820 $Y=21110 $D=111
M6566 474 2274 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=118220 $Y=21110 $D=111
M6567 VDD clk 2284 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=119330 $Y=45750 $D=111
M6568 2292 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=119730 $Y=45110 $D=111
M6569 2286 2289 2292 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=120130 $Y=45350 $D=111
M6570 VDD 2284 2289 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=121070 $Y=44790 $D=111
M6571 2285 475 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=121470 $Y=45590 $D=111
M6572 2293 2289 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=122390 $Y=44790 $D=111
M6573 2287 2285 2293 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=122710 $Y=44790 $D=111
M6574 2295 2286 2287 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=123240 $Y=45630 $D=111
M6575 VDD 2288 2295 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=123560 $Y=45630 $D=111
M6576 2288 2287 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=123960 $Y=45110 $D=111
M6577 VDD 2287 2288 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=124440 $Y=45110 $D=111
M6578 2288 543 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=124880 $Y=45510 $D=111
M6579 2291 2286 2288 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=125360 $Y=45170 $D=111
M6580 2288 2286 2291 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=125840 $Y=45110 $D=111
M6581 2300 2290 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=126700 $Y=45110 $D=111
M6582 2291 2289 2300 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=127020 $Y=45110 $D=111
M6583 VDD 543 2291 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=127500 $Y=44990 $D=111
M6584 VDD 2291 2290 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=127820 $Y=45810 $D=111
M6585 444 2291 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=128220 $Y=44790 $D=111
M6586 VDD clk 2301 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=134930 $Y=24150 $D=111
M6587 2309 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=135330 $Y=23510 $D=111
M6588 2303 2306 2309 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=135730 $Y=23750 $D=111
M6589 VDD 2301 2306 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=136670 $Y=23190 $D=111
M6590 2302 852 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=137070 $Y=23990 $D=111
M6591 2310 2306 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=137990 $Y=23190 $D=111
M6592 2304 2302 2310 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=138310 $Y=23190 $D=111
M6593 2312 2303 2304 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=138840 $Y=24030 $D=111
M6594 VDD 2305 2312 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=139160 $Y=24030 $D=111
M6595 2305 2304 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=139560 $Y=23510 $D=111
M6596 VDD 2304 2305 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=140040 $Y=23510 $D=111
M6597 2305 479 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=140480 $Y=23910 $D=111
M6598 2308 2303 2305 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=140960 $Y=23570 $D=111
M6599 2305 2303 2308 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=141440 $Y=23510 $D=111
M6600 2317 2307 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=142300 $Y=23510 $D=111
M6601 2308 2306 2317 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=142620 $Y=23510 $D=111
M6602 VDD 479 2308 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=143100 $Y=23390 $D=111
M6603 VDD 2308 2307 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=143420 $Y=24210 $D=111
M6604 505 2308 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=143820 $Y=23190 $D=111
M6605 VDD clk 2318 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=146130 $Y=71510 $D=111
M6606 2326 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=146530 $Y=71510 $D=111
M6607 2320 2323 2326 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=146930 $Y=71510 $D=111
M6608 VDD 2318 2323 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=147870 $Y=71650 $D=111
M6609 2319 552 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=148270 $Y=71650 $D=111
M6610 2327 2323 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=149190 $Y=71790 $D=111
M6611 2321 2319 2327 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=149510 $Y=71790 $D=111
M6612 2329 2320 2321 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=150040 $Y=71690 $D=111
M6613 VDD 2322 2329 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=150360 $Y=71690 $D=111
M6614 2322 2321 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=150760 $Y=71690 $D=111
M6615 VDD 2321 2322 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=151240 $Y=71690 $D=111
M6616 2322 610 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=151680 $Y=71690 $D=111
M6617 2325 2320 2322 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=152160 $Y=71690 $D=111
M6618 2322 2320 2325 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=152640 $Y=71690 $D=111
M6619 2334 2324 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=153500 $Y=72210 $D=111
M6620 2325 2323 2334 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=153820 $Y=72210 $D=111
M6621 VDD 610 2325 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=154300 $Y=72210 $D=111
M6622 VDD 2325 2324 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=154620 $Y=71510 $D=111
M6623 617 2325 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=155020 $Y=71510 $D=111
M6624 VDD clk 2335 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=149330 $Y=35510 $D=111
M6625 2343 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=149730 $Y=35510 $D=111
M6626 2337 2340 2343 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=150130 $Y=35510 $D=111
M6627 VDD 2335 2340 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=151070 $Y=35650 $D=111
M6628 2336 596 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=151470 $Y=35650 $D=111
M6629 2344 2340 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=152390 $Y=35790 $D=111
M6630 2338 2336 2344 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=152710 $Y=35790 $D=111
M6631 2346 2337 2338 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=153240 $Y=35690 $D=111
M6632 VDD 2339 2346 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=153560 $Y=35690 $D=111
M6633 2339 2338 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=153960 $Y=35690 $D=111
M6634 VDD 2338 2339 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=154440 $Y=35690 $D=111
M6635 2339 564 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=154880 $Y=35690 $D=111
M6636 2342 2337 2339 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=155360 $Y=35690 $D=111
M6637 2339 2337 2342 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=155840 $Y=35690 $D=111
M6638 2351 2341 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=156700 $Y=36210 $D=111
M6639 2342 2340 2351 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=157020 $Y=36210 $D=111
M6640 VDD 564 2342 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=157500 $Y=36210 $D=111
M6641 VDD 2342 2341 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=157820 $Y=35510 $D=111
M6642 632 2342 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=158220 $Y=35510 $D=111
M6643 VDD clk 2352 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=150530 $Y=45750 $D=111
M6644 2360 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=150930 $Y=45110 $D=111
M6645 2354 2357 2360 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=151330 $Y=45350 $D=111
M6646 VDD 2352 2357 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=152270 $Y=44790 $D=111
M6647 2353 606 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=152670 $Y=45590 $D=111
M6648 2361 2357 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=153590 $Y=44790 $D=111
M6649 2355 2353 2361 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=153910 $Y=44790 $D=111
M6650 2363 2354 2355 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=154440 $Y=45630 $D=111
M6651 VDD 2356 2363 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=154760 $Y=45630 $D=111
M6652 2356 2355 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=155160 $Y=45110 $D=111
M6653 VDD 2355 2356 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=155640 $Y=45110 $D=111
M6654 2356 697 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=156080 $Y=45510 $D=111
M6655 2359 2354 2356 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=156560 $Y=45170 $D=111
M6656 2356 2354 2359 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=157040 $Y=45110 $D=111
M6657 2368 2358 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=157900 $Y=45110 $D=111
M6658 2359 2357 2368 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=158220 $Y=45110 $D=111
M6659 VDD 697 2359 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=158700 $Y=44990 $D=111
M6660 VDD 2359 2358 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=159020 $Y=45810 $D=111
M6661 646 2359 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=159420 $Y=44790 $D=111
M6662 VDD clk 2369 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=156530 $Y=64310 $D=111
M6663 2377 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=156930 $Y=64310 $D=111
M6664 2371 2374 2377 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=157330 $Y=64310 $D=111
M6665 VDD 2369 2374 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=158270 $Y=64450 $D=111
M6666 2370 858 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=158670 $Y=64450 $D=111
M6667 2378 2374 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=159590 $Y=64590 $D=111
M6668 2372 2370 2378 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=159910 $Y=64590 $D=111
M6669 2380 2371 2372 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=160440 $Y=64490 $D=111
M6670 VDD 2373 2380 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=160760 $Y=64490 $D=111
M6671 2373 2372 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=161160 $Y=64490 $D=111
M6672 VDD 2372 2373 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=161640 $Y=64490 $D=111
M6673 2373 610 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=162080 $Y=64490 $D=111
M6674 2376 2371 2373 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=162560 $Y=64490 $D=111
M6675 2373 2371 2376 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=163040 $Y=64490 $D=111
M6676 2385 2375 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=163900 $Y=65010 $D=111
M6677 2376 2374 2385 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=164220 $Y=65010 $D=111
M6678 VDD 610 2376 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=164700 $Y=65010 $D=111
M6679 VDD 2376 2375 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=165020 $Y=64310 $D=111
M6680 652 2376 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=165420 $Y=64310 $D=111
M6681 VDD clk 2386 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=159330 $Y=35510 $D=111
M6682 2394 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=159730 $Y=35510 $D=111
M6683 2388 2391 2394 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=160130 $Y=35510 $D=111
M6684 VDD 2386 2391 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=161070 $Y=35650 $D=111
M6685 2387 694 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=161470 $Y=35650 $D=111
M6686 2395 2391 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=162390 $Y=35790 $D=111
M6687 2389 2387 2395 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=162710 $Y=35790 $D=111
M6688 2397 2388 2389 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=163240 $Y=35690 $D=111
M6689 VDD 2390 2397 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=163560 $Y=35690 $D=111
M6690 2390 2389 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=163960 $Y=35690 $D=111
M6691 VDD 2389 2390 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=164440 $Y=35690 $D=111
M6692 2390 760 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=164880 $Y=35690 $D=111
M6693 2393 2388 2390 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=165360 $Y=35690 $D=111
M6694 2390 2388 2393 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=165840 $Y=35690 $D=111
M6695 2402 2392 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=166700 $Y=36210 $D=111
M6696 2393 2391 2402 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=167020 $Y=36210 $D=111
M6697 VDD 760 2393 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=167500 $Y=36210 $D=111
M6698 VDD 2393 2392 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=167820 $Y=35510 $D=111
M6699 683 2393 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=168220 $Y=35510 $D=111
M6700 VDD clk 2403 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=164130 $Y=71510 $D=111
M6701 2411 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=164530 $Y=71510 $D=111
M6702 2405 2408 2411 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=164930 $Y=71510 $D=111
M6703 VDD 2403 2408 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=165870 $Y=71650 $D=111
M6704 2404 859 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=166270 $Y=71650 $D=111
M6705 2412 2408 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=167190 $Y=71790 $D=111
M6706 2406 2404 2412 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=167510 $Y=71790 $D=111
M6707 2414 2405 2406 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=168040 $Y=71690 $D=111
M6708 VDD 2407 2414 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=168360 $Y=71690 $D=111
M6709 2407 2406 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=168760 $Y=71690 $D=111
M6710 VDD 2406 2407 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=169240 $Y=71690 $D=111
M6711 2407 610 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=169680 $Y=71690 $D=111
M6712 2410 2405 2407 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=170160 $Y=71690 $D=111
M6713 2407 2405 2410 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=170640 $Y=71690 $D=111
M6714 2419 2409 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=171500 $Y=72210 $D=111
M6715 2410 2408 2419 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=171820 $Y=72210 $D=111
M6716 VDD 610 2410 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=172300 $Y=72210 $D=111
M6717 VDD 2410 2409 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=172620 $Y=71510 $D=111
M6718 576 2410 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=173020 $Y=71510 $D=111
M6719 VDD clk 2420 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=169730 $Y=28310 $D=111
M6720 2428 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=170130 $Y=28310 $D=111
M6721 2422 2425 2428 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=170530 $Y=28310 $D=111
M6722 VDD 2420 2425 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=171470 $Y=28450 $D=111
M6723 2421 704 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=171870 $Y=28450 $D=111
M6724 2429 2425 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=172790 $Y=28590 $D=111
M6725 2423 2421 2429 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=173110 $Y=28590 $D=111
M6726 2431 2422 2423 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=173640 $Y=28490 $D=111
M6727 VDD 2424 2431 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=173960 $Y=28490 $D=111
M6728 2424 2423 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=174360 $Y=28490 $D=111
M6729 VDD 2423 2424 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=174840 $Y=28490 $D=111
M6730 2424 706 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=175280 $Y=28490 $D=111
M6731 2427 2422 2424 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=175760 $Y=28490 $D=111
M6732 2424 2422 2427 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=176240 $Y=28490 $D=111
M6733 2436 2426 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=177100 $Y=29010 $D=111
M6734 2427 2425 2436 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=177420 $Y=29010 $D=111
M6735 VDD 706 2427 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=177900 $Y=29010 $D=111
M6736 VDD 2427 2426 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=178220 $Y=28310 $D=111
M6737 716 2427 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=178620 $Y=28310 $D=111
M6738 VDD clk 2437 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=175730 $Y=13910 $D=111
M6739 2445 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=176130 $Y=13910 $D=111
M6740 2439 2442 2445 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=176530 $Y=13910 $D=111
M6741 VDD 2437 2442 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=177470 $Y=14050 $D=111
M6742 2438 754 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=177870 $Y=14050 $D=111
M6743 2446 2442 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=178790 $Y=14190 $D=111
M6744 2440 2438 2446 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=179110 $Y=14190 $D=111
M6745 2448 2439 2440 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=179640 $Y=14090 $D=111
M6746 VDD 2441 2448 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=179960 $Y=14090 $D=111
M6747 2441 2440 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=180360 $Y=14090 $D=111
M6748 VDD 2440 2441 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=180840 $Y=14090 $D=111
M6749 2441 706 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=181280 $Y=14090 $D=111
M6750 2444 2439 2441 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=181760 $Y=14090 $D=111
M6751 2441 2439 2444 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=182240 $Y=14090 $D=111
M6752 2453 2443 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=183100 $Y=14610 $D=111
M6753 2444 2442 2453 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=183420 $Y=14610 $D=111
M6754 VDD 706 2444 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=183900 $Y=14610 $D=111
M6755 VDD 2444 2443 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=184220 $Y=13910 $D=111
M6756 733 2444 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=184620 $Y=13910 $D=111
M6757 VDD clk 2454 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=175730 $Y=67350 $D=111
M6758 2462 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=176130 $Y=66710 $D=111
M6759 2456 2459 2462 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=176530 $Y=66950 $D=111
M6760 VDD 2454 2459 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=177470 $Y=66390 $D=111
M6761 2455 762 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=177870 $Y=67190 $D=111
M6762 2463 2459 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=178790 $Y=66390 $D=111
M6763 2457 2455 2463 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=179110 $Y=66390 $D=111
M6764 2465 2456 2457 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=179640 $Y=67230 $D=111
M6765 VDD 2458 2465 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=179960 $Y=67230 $D=111
M6766 2458 2457 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=180360 $Y=66710 $D=111
M6767 VDD 2457 2458 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=180840 $Y=66710 $D=111
M6768 2458 760 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=181280 $Y=67110 $D=111
M6769 2461 2456 2458 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=181760 $Y=66770 $D=111
M6770 2458 2456 2461 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=182240 $Y=66710 $D=111
M6771 2470 2460 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=183100 $Y=66710 $D=111
M6772 2461 2459 2470 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=183420 $Y=66710 $D=111
M6773 VDD 760 2461 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=183900 $Y=66590 $D=111
M6774 VDD 2461 2460 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=184220 $Y=67410 $D=111
M6775 746 2461 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=184620 $Y=66390 $D=111
M6776 VDD clk 2471 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=176130 $Y=35510 $D=111
M6777 2479 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=176530 $Y=35510 $D=111
M6778 2473 2476 2479 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=176930 $Y=35510 $D=111
M6779 VDD 2471 2476 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=177870 $Y=35650 $D=111
M6780 2472 782 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=178270 $Y=35650 $D=111
M6781 2480 2476 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=179190 $Y=35790 $D=111
M6782 2474 2472 2480 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=179510 $Y=35790 $D=111
M6783 2482 2473 2474 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=180040 $Y=35690 $D=111
M6784 VDD 2475 2482 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=180360 $Y=35690 $D=111
M6785 2475 2474 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=180760 $Y=35690 $D=111
M6786 VDD 2474 2475 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=181240 $Y=35690 $D=111
M6787 2475 706 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=181680 $Y=35690 $D=111
M6788 2478 2473 2475 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=182160 $Y=35690 $D=111
M6789 2475 2473 2478 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=182640 $Y=35690 $D=111
M6790 2487 2477 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=183500 $Y=36210 $D=111
M6791 2478 2476 2487 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=183820 $Y=36210 $D=111
M6792 VDD 706 2478 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=184300 $Y=36210 $D=111
M6793 VDD 2478 2477 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=184620 $Y=35510 $D=111
M6794 717 2478 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=185020 $Y=35510 $D=111
M6795 VDD clk 2488 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07846e-13 as=1.088e-13 pd=8.43041e-07 ps=1.32e-06 nrd=0.932921 nrs=0.941176 sa=3.2e-07 sb=1.12e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=4.8e-15 panw8=0 panw9=0 panw10=0 $X=177730 $Y=49910 $D=111
M6796 2496 clk VDD VDD lppfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.45405e-13 as=3.10849e-13 pd=1.43581e-06 ps=2.42994e-06 nrd=0.1514 nrs=0.323666 sa=4.71327e-07 sb=5.92653e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=178130 $Y=49910 $D=111
M6797 2490 2493 2496 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.368e-13 as=1.09795e-13 pd=2.12e-06 ps=1.08419e-06 nrd=0.432432 nrs=0.200503 sa=8.71757e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-15 panw10=0 $X=178530 $Y=49910 $D=111
M6798 VDD 2488 2493 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.74945e-13 as=2.656e-13 pd=2.93702e-06 ps=2.96e-06 nrd=0.204329 nrs=0.197384 sa=2.28966e-07 sb=5.95862e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=179470 $Y=50050 $D=111
M6799 2489 864 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.056e-13 as=8.53277e-14 pd=1.36e-06 ps=9.11489e-07 nrd=0.814815 nrs=0.658392 sa=6.93333e-07 sb=2.93333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.2e-15 panw8=0 panw9=0 panw10=0 $X=179870 $Y=50050 $D=111
M6800 2497 2493 VDD VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02e-13 as=2.41762e-13 pd=1.22e-06 ps=2.58255e-06 nrd=0.0980392 nrs=0.232374 sa=4.07059e-07 sb=8.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=180790 $Y=50190 $D=111
M6801 2491 2489 2497 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.84502e-13 as=1.02e-13 pd=2.40092e-06 ps=1.22e-06 nrd=0.273454 nrs=0.0980392 sa=7.27059e-07 sb=6.16471e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=181110 $Y=50190 $D=111
M6802 2499 2490 2491 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=7.80985e-14 pd=4.8e-07 ps=6.59077e-07 nrd=0.357143 nrs=0.996154 sa=7.46429e-07 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=181640 $Y=50090 $D=111
M6803 VDD 2492 2499 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.55176e-14 as=2.8e-14 pd=7.53529e-07 ps=4.8e-07 nrd=0.963235 nrs=0.357143 sa=1.06643e-06 sb=2e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=181960 $Y=50090 $D=111
M6804 2492 2491 VDD VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.44e-13 as=2.15765e-13 pd=1.16e-06 ps=2.15294e-06 nrd=0.225 nrs=0.337132 sa=6.6725e-07 sb=1.36e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=182360 $Y=50090 $D=111
M6805 VDD 2491 2492 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9027e-13 as=1.44e-13 pd=1.97838e-06 ps=1.16e-06 nrd=0.297297 nrs=0.225 sa=1.091e-06 sb=9.62e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=182840 $Y=50090 $D=111
M6806 2492 760 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.4386e-14 as=9.51351e-14 pd=7.7193e-07 ps=9.89189e-07 nrd=0.464912 nrs=0.594595 sa=1.696e-06 sb=1.244e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=183280 $Y=50090 $D=111
M6807 2495 2490 2492 VDD lppfet w=7.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.33777e-13 as=1.37614e-13 pd=1.11481e-06 ps=1.42807e-06 nrd=0.244296 nrs=0.251304 sa=1.10811e-06 sb=7.25405e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=183760 $Y=50090 $D=111
M6808 2492 2490 2495 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.936e-13 as=1.44623e-13 pd=2.24e-06 ps=1.20519e-06 nrd=0.3025 nrs=0.225974 sa=1.304e-06 sb=2.42e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=184240 $Y=50090 $D=111
M6809 2504 2494 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.512e-13 pd=4.8e-07 ps=1.64e-06 nrd=0.357143 nrs=1.92857 sa=3.6e-07 sb=1.87e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.68e-14 panw9=1.68e-14 panw10=0 $X=185100 $Y=50610 $D=111
M6810 2495 2493 2504 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.53412e-14 as=2.8e-14 pd=6.25882e-07 ps=4.8e-07 nrd=0.705882 nrs=0.357143 sa=6.8e-07 sb=1.55e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.26e-14 panw9=2.1e-14 panw10=0 $X=185420 $Y=50610 $D=111
M6811 VDD 760 2495 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02303e-13 as=7.90588e-14 pd=8e-07 ps=8.94118e-07 nrd=0.639394 nrs=0.494118 sa=8.96e-07 sb=1.07e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=4.8e-14 panw10=0 $X=185900 $Y=50610 $D=111
M6812 VDD 2495 2494 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.16121e-14 as=1.008e-13 pd=5.6e-07 ps=1.28e-06 nrd=0.91342 nrs=1.28571 sa=3.6e-07 sb=7.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=186220 $Y=49910 $D=111
M6813 726 2495 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.55e-13 as=3.32485e-13 pd=3.3e-06 ps=2.6e-06 nrd=0.269231 nrs=0.196737 sa=8.05538e-07 sb=3.5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=186620 $Y=49910 $D=111
M6814 VDD 256 2505 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=69930 $Y=13910 $D=111
M6815 2505 264 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=70390 $Y=13910 $D=111
M6816 2506 310 2505 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=70880 $Y=13910 $D=111
M6817 VDD 2506 251 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=6.87619e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=71350 $Y=15040 $D=111
M6818 2505 result[1] 2506 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=71360 $Y=13910 $D=111
M6819 VDD 256 2509 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=76330 $Y=13910 $D=111
M6820 2509 143 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=76790 $Y=13910 $D=111
M6821 2510 310 2509 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=77280 $Y=13910 $D=111
M6822 VDD 2510 828 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=5.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=77750 $Y=15040 $D=111
M6823 2509 result[2] 2510 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=77760 $Y=13910 $D=111
M6824 VDD 256 2513 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=79130 $Y=13910 $D=111
M6825 2513 298 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=79590 $Y=13910 $D=111
M6826 2514 310 2513 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=80080 $Y=13910 $D=111
M6827 VDD 2514 269 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=5.61429e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=80550 $Y=15040 $D=111
M6828 2513 result[0] 2514 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=80560 $Y=13910 $D=111
M6829 VDD 300 2517 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=79930 $Y=31390 $D=111
M6830 2517 159 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=80390 $Y=31390 $D=111
M6831 2518 306 2517 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=80880 $Y=31390 $D=111
M6832 305 2518 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=1.29429e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=81350 $Y=30440 $D=111
M6833 2517 result[5] 2518 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=81360 $Y=31390 $D=111
M6834 VDD 300 2521 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=82730 $Y=31390 $D=111
M6835 2521 109 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=83190 $Y=31390 $D=111
M6836 2522 306 2521 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=83680 $Y=31390 $D=111
M6837 321 2522 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=5.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=84150 $Y=30440 $D=111
M6838 2521 result[6] 2522 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=84160 $Y=31390 $D=111
M6839 VDD 318 2525 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=85530 $Y=21110 $D=111
M6840 2525 62 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=85990 $Y=21110 $D=111
M6841 2526 345 2525 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=86480 $Y=21110 $D=111
M6842 VDD 2526 322 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=5.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=86950 $Y=22240 $D=111
M6843 2525 result[4] 2526 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=86960 $Y=21110 $D=111
M6844 VDD 389 2529 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=88330 $Y=13910 $D=111
M6845 2529 100 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=88790 $Y=13910 $D=111
M6846 2530 326 2529 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=89280 $Y=13910 $D=111
M6847 VDD 2530 333 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=1.51857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=89750 $Y=15040 $D=111
M6848 2529 result[3] 2530 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=89760 $Y=13910 $D=111
M6849 VDD 318 2533 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=88730 $Y=21110 $D=111
M6850 2533 260 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=89190 $Y=21110 $D=111
M6851 2534 345 2533 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=89680 $Y=21110 $D=111
M6852 VDD 2534 332 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=7.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=90150 $Y=22240 $D=111
M6853 2533 result[7] 2534 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=90160 $Y=21110 $D=111
M6854 VDD 377 2537 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=95930 $Y=21110 $D=111
M6855 2537 239 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=96390 $Y=21110 $D=111
M6856 2538 368 2537 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=96880 $Y=21110 $D=111
M6857 VDD 2538 832 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=1.51857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=97350 $Y=22240 $D=111
M6858 2537 result[8] 2538 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=97360 $Y=21110 $D=111
M6859 VDD 389 2541 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=97130 $Y=13910 $D=111
M6860 2541 359 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=97590 $Y=13910 $D=111
M6861 2542 326 2541 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=98080 $Y=13910 $D=111
M6862 VDD 2542 364 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=5.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=98550 $Y=15040 $D=111
M6863 2541 result[10] 2542 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=98560 $Y=13910 $D=111
M6864 VDD 399 2545 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=99930 $Y=21110 $D=111
M6865 2545 363 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=100390 $Y=21110 $D=111
M6866 2546 368 2545 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=100880 $Y=21110 $D=111
M6867 VDD 2546 373 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=5.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=101350 $Y=22240 $D=111
M6868 2545 result[9] 2546 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=101360 $Y=21110 $D=111
M6869 VDD 389 2549 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=102330 $Y=13910 $D=111
M6870 2549 418 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=102790 $Y=13910 $D=111
M6871 2550 326 2549 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=103280 $Y=13910 $D=111
M6872 VDD 2550 385 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=1.51857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=103750 $Y=15040 $D=111
M6873 2549 result[11] 2550 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=103760 $Y=13910 $D=111
M6874 VDD 408 2553 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=106730 $Y=16990 $D=111
M6875 2553 452 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=107190 $Y=16990 $D=111
M6876 2554 396 2553 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=107680 $Y=16990 $D=111
M6877 388 2554 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=5.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=108150 $Y=16040 $D=111
M6878 2553 result[12] 2554 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=108160 $Y=16990 $D=111
M6879 VDD 408 2557 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=118730 $Y=16990 $D=111
M6880 2557 444 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=119190 $Y=16990 $D=111
M6881 2558 396 2557 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=119680 $Y=16990 $D=111
M6882 453 2558 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=5.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=120150 $Y=16040 $D=111
M6883 2557 result[14] 2558 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=120160 $Y=16990 $D=111
M6884 VDD 408 2561 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=118730 $Y=24190 $D=111
M6885 2561 839 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=119190 $Y=24190 $D=111
M6886 2562 396 2561 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=119680 $Y=24190 $D=111
M6887 454 2562 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=7.24286e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=120150 $Y=23240 $D=111
M6888 2561 result[13] 2562 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=120160 $Y=24190 $D=111
M6889 VDD 491 2565 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=123530 $Y=13910 $D=111
M6890 2565 456 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=123990 $Y=13910 $D=111
M6891 2566 526 2565 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=124480 $Y=13910 $D=111
M6892 VDD 2566 424 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=6.93333e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=124950 $Y=15040 $D=111
M6893 2565 result[15] 2566 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=124960 $Y=13910 $D=111
M6894 VDD 491 2569 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=126330 $Y=13910 $D=111
M6895 2569 474 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=126790 $Y=13910 $D=111
M6896 2570 526 2569 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=127280 $Y=13910 $D=111
M6897 VDD 2570 449 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=127750 $Y=15040 $D=111
M6898 2569 result[16] 2570 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=127760 $Y=13910 $D=111
M6899 VDD 500 2573 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=131130 $Y=13910 $D=111
M6900 2573 505 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=131590 $Y=13910 $D=111
M6901 2574 526 2573 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=132080 $Y=13910 $D=111
M6902 VDD 2574 513 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=132550 $Y=15040 $D=111
M6903 2573 result[17] 2574 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=132560 $Y=13910 $D=111
M6904 VDD 500 2577 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=136730 $Y=13910 $D=111
M6905 2577 568 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=137190 $Y=13910 $D=111
M6906 2578 570 2577 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=137680 $Y=13910 $D=111
M6907 VDD 2578 541 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=138150 $Y=15040 $D=111
M6908 2577 result[18] 2578 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=138160 $Y=13910 $D=111
M6909 VDD 611 2581 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=145130 $Y=16990 $D=111
M6910 2581 632 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=145590 $Y=16990 $D=111
M6911 2582 570 2581 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=146080 $Y=16990 $D=111
M6912 579 2582 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=5.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=146550 $Y=16040 $D=111
M6913 2581 result[19] 2582 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=146560 $Y=16990 $D=111
M6914 VDD 593 2585 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=150330 $Y=16990 $D=111
M6915 2585 597 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=150790 $Y=16990 $D=111
M6916 2586 620 2585 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=151280 $Y=16990 $D=111
M6917 604 2586 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=7.31429e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=151750 $Y=16040 $D=111
M6918 2585 result[21] 2586 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=151760 $Y=16990 $D=111
M6919 VDD 593 2589 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=154730 $Y=16990 $D=111
M6920 2589 646 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=155190 $Y=16990 $D=111
M6921 2590 570 2589 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=155680 $Y=16990 $D=111
M6922 623 2590 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=5.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=156150 $Y=16040 $D=111
M6923 2589 result[20] 2590 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=156160 $Y=16990 $D=111
M6924 VDD 688 2593 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=156330 $Y=31390 $D=111
M6925 2593 652 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=156790 $Y=31390 $D=111
M6926 2594 651 2593 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=157280 $Y=31390 $D=111
M6927 612 2594 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=6.87619e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=157750 $Y=30440 $D=111
M6928 2593 result[25] 2594 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=157760 $Y=31390 $D=111
M6929 VDD 593 2597 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=157530 $Y=16990 $D=111
M6930 2597 609 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=157990 $Y=16990 $D=111
M6931 2598 645 2597 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=158480 $Y=16990 $D=111
M6932 621 2598 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=6.74762e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=158950 $Y=16040 $D=111
M6933 2597 result[22] 2598 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=158960 $Y=16990 $D=111
M6934 VDD 682 2601 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=157530 $Y=24190 $D=111
M6935 2601 576 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=157990 $Y=24190 $D=111
M6936 2602 620 2601 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=158480 $Y=24190 $D=111
M6937 563 2602 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=6.87619e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=158950 $Y=23240 $D=111
M6938 2601 result[24] 2602 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=158960 $Y=24190 $D=111
M6939 VDD 682 2605 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=160330 $Y=24190 $D=111
M6940 2605 617 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=160790 $Y=24190 $D=111
M6941 2606 620 2605 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=161280 $Y=24190 $D=111
M6942 654 2606 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=5.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=161750 $Y=23240 $D=111
M6943 2605 result[23] 2606 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=161760 $Y=24190 $D=111
M6944 VDD 689 2609 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=161530 $Y=31390 $D=111
M6945 2609 746 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=161990 $Y=31390 $D=111
M6946 2610 651 2609 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=162480 $Y=31390 $D=111
M6947 656 2610 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=5.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=162950 $Y=30440 $D=111
M6948 2609 result[26] 2610 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=162960 $Y=31390 $D=111
M6949 VDD 688 2613 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=164730 $Y=16990 $D=111
M6950 2613 683 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=165190 $Y=16990 $D=111
M6951 2614 701 2613 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=165680 $Y=16990 $D=111
M6952 643 2614 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=9.94762e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=166150 $Y=16040 $D=111
M6953 2613 result[28] 2614 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=166160 $Y=16990 $D=111
M6954 VDD 682 2617 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=166330 $Y=24190 $D=111
M6955 2617 726 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=166790 $Y=24190 $D=111
M6956 2618 651 2617 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=167280 $Y=24190 $D=111
M6957 678 2618 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=6.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=167750 $Y=23240 $D=111
M6958 2617 result[27] 2618 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=167760 $Y=24190 $D=111
M6959 VDD 688 2621 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=169930 $Y=13910 $D=111
M6960 2621 717 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=170390 $Y=13910 $D=111
M6961 2622 701 2621 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=170880 $Y=13910 $D=111
M6962 VDD 2622 699 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=5.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=171350 $Y=15040 $D=111
M6963 2621 result[29] 2622 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=171360 $Y=13910 $D=111
M6964 VDD 693 2625 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=172730 $Y=13910 $D=111
M6965 2625 716 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=173190 $Y=13910 $D=111
M6966 2626 701 2625 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=173680 $Y=13910 $D=111
M6967 VDD 2626 708 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.72e-14 as=1.344e-13 pd=7.4e-07 ps=1.48e-06 nrd=0.380952 nrs=0.761905 sa=3.2e-07 sb=5.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=174150 $Y=15040 $D=111
M6968 2625 result[30] 2626 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=174160 $Y=13910 $D=111
M6969 VDD 693 2629 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41682e-13 as=2e-13 pd=1.38409e-06 ps=2.5e-06 nrd=1.57424 nrs=2.22222 sa=2.4e-07 sb=1.75e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=177130 $Y=16990 $D=111
M6970 2629 733 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.55e-14 as=1.41682e-13 pd=6.7e-07 ps=1.38409e-06 nrd=0.616667 nrs=1.57424 sa=7e-07 sb=1.29e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=177590 $Y=16990 $D=111
M6971 2630 701 2629 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.4e-14 as=5.55e-14 pd=6.6e-07 ps=6.7e-07 nrd=0.6 nrs=0.616667 sa=1.19e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=178080 $Y=16990 $D=111
M6972 740 2630 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.344e-13 as=6.72e-14 pd=1.48e-06 ps=7.4e-07 nrd=0.761905 nrs=0.380952 sa=5.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=5.04e-14 $X=178550 $Y=16040 $D=111
M6973 2629 result[31] 2630 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=5.4e-14 pd=1.24e-06 ps=6.6e-07 nrd=1.06667 nrs=0.6 sa=1.67e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=178560 $Y=16990 $D=111
M6974 2641 78 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=25660 $Y=14640 $D=111
M6975 2634 2636 2641 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=25980 $Y=14640 $D=111
M6976 VDD 68 2634 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=26460 $Y=14640 $D=111
M6977 VDD clk 2633 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=26980 $Y=13910 $D=111
M6978 2636 2633 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=27490 $Y=13950 $D=111
M6979 2643 2633 2634 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=28050 $Y=14410 $D=111
M6980 VDD 2635 2643 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=28370 $Y=14410 $D=111
M6981 2635 2634 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=28910 $Y=14410 $D=111
M6982 2637 2633 2635 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=29740 $Y=14660 $D=111
M6983 2646 2636 2637 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=30470 $Y=14660 $D=111
M6984 VDD 2639 2646 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=30800 $Y=14660 $D=111
M6985 2639 68 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=31260 $Y=14590 $D=111
M6986 VDD 2637 2639 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=31820 $Y=14880 $D=111
M6987 2638 2639 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=32430 $Y=14240 $D=111
M6988 VDD 2638 919 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=33370 $Y=14050 $D=111
M6989 weight_out[3] 2639 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=33870 $Y=14050 $D=111
M6990 2657 269 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=72060 $Y=16280 $D=111
M6991 2650 2652 2657 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=72380 $Y=16280 $D=111
M6992 VDD 316 2650 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=72860 $Y=16280 $D=111
M6993 VDD clk 2649 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=73380 $Y=16870 $D=111
M6994 2652 2649 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=73890 $Y=16970 $D=111
M6995 2659 2649 2650 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=74450 $Y=16510 $D=111
M6996 VDD 2651 2659 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=74770 $Y=16510 $D=111
M6997 2651 2650 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=75310 $Y=16510 $D=111
M6998 2653 2649 2651 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=76140 $Y=16260 $D=111
M6999 2662 2652 2653 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=76870 $Y=16260 $D=111
M7000 VDD 2655 2662 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=77200 $Y=16260 $D=111
M7001 2655 316 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=77660 $Y=16330 $D=111
M7002 VDD 2653 2655 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=78220 $Y=16040 $D=111
M7003 2654 2655 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=78830 $Y=16680 $D=111
M7004 VDD 2654 920 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=79770 $Y=16810 $D=111
M7005 result[0] 2655 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=80270 $Y=16810 $D=111
M7006 2673 322 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=82060 $Y=16280 $D=111
M7007 2666 2668 2673 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=82380 $Y=16280 $D=111
M7008 VDD 316 2666 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=82860 $Y=16280 $D=111
M7009 VDD clk 2665 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=83380 $Y=16870 $D=111
M7010 2668 2665 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=83890 $Y=16970 $D=111
M7011 2675 2665 2666 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=84450 $Y=16510 $D=111
M7012 VDD 2667 2675 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=84770 $Y=16510 $D=111
M7013 2667 2666 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=85310 $Y=16510 $D=111
M7014 2669 2665 2667 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=86140 $Y=16260 $D=111
M7015 2678 2668 2669 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=86870 $Y=16260 $D=111
M7016 VDD 2671 2678 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=87200 $Y=16260 $D=111
M7017 2671 316 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=87660 $Y=16330 $D=111
M7018 VDD 2669 2671 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=88220 $Y=16040 $D=111
M7019 2670 2671 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=88830 $Y=16680 $D=111
M7020 VDD 2670 921 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=89770 $Y=16810 $D=111
M7021 result[4] 2671 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=90270 $Y=16810 $D=111
M7022 2689 321 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=87260 $Y=30680 $D=111
M7023 2682 2684 2689 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=87580 $Y=30680 $D=111
M7024 VDD 303 2682 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=88060 $Y=30680 $D=111
M7025 VDD clk 2681 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=88580 $Y=31270 $D=111
M7026 2684 2681 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=89090 $Y=31370 $D=111
M7027 2691 2681 2682 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=89650 $Y=30910 $D=111
M7028 VDD 2683 2691 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=89970 $Y=30910 $D=111
M7029 2683 2682 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=90510 $Y=30910 $D=111
M7030 2685 2681 2683 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=91340 $Y=30660 $D=111
M7031 2694 2684 2685 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=92070 $Y=30660 $D=111
M7032 VDD 2687 2694 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=92400 $Y=30660 $D=111
M7033 2687 303 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=92860 $Y=30730 $D=111
M7034 VDD 2685 2687 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=93420 $Y=30440 $D=111
M7035 2686 2687 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=94030 $Y=31080 $D=111
M7036 VDD 2686 922 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=94970 $Y=31210 $D=111
M7037 result[6] 2687 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=95470 $Y=31210 $D=111
M7038 2705 192 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=95660 $Y=36240 $D=111
M7039 2698 2700 2705 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=95980 $Y=36240 $D=111
M7040 VDD 374 2698 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=96460 $Y=36240 $D=111
M7041 VDD clk 2697 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=96980 $Y=35510 $D=111
M7042 2700 2697 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=97490 $Y=35550 $D=111
M7043 2707 2697 2698 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=98050 $Y=36010 $D=111
M7044 VDD 2699 2707 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=98370 $Y=36010 $D=111
M7045 2699 2698 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=98910 $Y=36010 $D=111
M7046 2701 2697 2699 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=99740 $Y=36260 $D=111
M7047 2710 2700 2701 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=100470 $Y=36260 $D=111
M7048 VDD 2703 2710 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=100800 $Y=36260 $D=111
M7049 2703 374 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=101260 $Y=36190 $D=111
M7050 VDD 2701 2703 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=101820 $Y=36480 $D=111
M7051 2702 2703 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=102430 $Y=35840 $D=111
M7052 VDD 2702 923 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=103370 $Y=35650 $D=111
M7053 data_out[3] 2703 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=103870 $Y=35650 $D=111
M7054 2721 373 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=96060 $Y=16280 $D=111
M7055 2714 2716 2721 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=96380 $Y=16280 $D=111
M7056 VDD 371 2714 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=96860 $Y=16280 $D=111
M7057 VDD clk 2713 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=97380 $Y=16870 $D=111
M7058 2716 2713 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=97890 $Y=16970 $D=111
M7059 2723 2713 2714 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=98450 $Y=16510 $D=111
M7060 VDD 2715 2723 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=98770 $Y=16510 $D=111
M7061 2715 2714 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=99310 $Y=16510 $D=111
M7062 2717 2713 2715 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=100140 $Y=16260 $D=111
M7063 2726 2716 2717 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=100870 $Y=16260 $D=111
M7064 VDD 2719 2726 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=101200 $Y=16260 $D=111
M7065 2719 371 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=101660 $Y=16330 $D=111
M7066 VDD 2717 2719 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=102220 $Y=16040 $D=111
M7067 2718 2719 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=102830 $Y=16680 $D=111
M7068 VDD 2718 924 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=103770 $Y=16810 $D=111
M7069 result[9] 2719 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=104270 $Y=16810 $D=111
M7070 2737 254 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=101660 $Y=29040 $D=111
M7071 2730 2732 2737 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=101980 $Y=29040 $D=111
M7072 VDD 374 2730 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=102460 $Y=29040 $D=111
M7073 VDD clk 2729 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=102980 $Y=28310 $D=111
M7074 2732 2729 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=103490 $Y=28350 $D=111
M7075 2739 2729 2730 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=104050 $Y=28810 $D=111
M7076 VDD 2731 2739 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=104370 $Y=28810 $D=111
M7077 2731 2730 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=104910 $Y=28810 $D=111
M7078 2733 2729 2731 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=105740 $Y=29060 $D=111
M7079 2742 2732 2733 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=106470 $Y=29060 $D=111
M7080 VDD 2735 2742 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=106800 $Y=29060 $D=111
M7081 2735 374 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=107260 $Y=28990 $D=111
M7082 VDD 2733 2735 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=107820 $Y=29280 $D=111
M7083 2734 2735 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=108430 $Y=28640 $D=111
M7084 VDD 2734 925 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=109370 $Y=28450 $D=111
M7085 data_out[2] 2735 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=109870 $Y=28450 $D=111
M7086 2753 385 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=105660 $Y=9080 $D=111
M7087 2746 2748 2753 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=105980 $Y=9080 $D=111
M7088 VDD 371 2746 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=106460 $Y=9080 $D=111
M7089 VDD clk 2745 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=106980 $Y=9670 $D=111
M7090 2748 2745 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=107490 $Y=9770 $D=111
M7091 2755 2745 2746 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=108050 $Y=9310 $D=111
M7092 VDD 2747 2755 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=108370 $Y=9310 $D=111
M7093 2747 2746 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=108910 $Y=9310 $D=111
M7094 2749 2745 2747 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=109740 $Y=9060 $D=111
M7095 2758 2748 2749 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=110470 $Y=9060 $D=111
M7096 VDD 2751 2758 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=110800 $Y=9060 $D=111
M7097 2751 371 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=111260 $Y=9130 $D=111
M7098 VDD 2749 2751 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=111820 $Y=8840 $D=111
M7099 2750 2751 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=112430 $Y=9480 $D=111
M7100 VDD 2750 926 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=113370 $Y=9610 $D=111
M7101 result[11] 2751 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=113870 $Y=9610 $D=111
M7102 2769 454 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=109660 $Y=16280 $D=111
M7103 2762 2764 2769 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=109980 $Y=16280 $D=111
M7104 VDD 428 2762 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=110460 $Y=16280 $D=111
M7105 VDD clk 2761 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=110980 $Y=16870 $D=111
M7106 2764 2761 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=111490 $Y=16970 $D=111
M7107 2771 2761 2762 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=112050 $Y=16510 $D=111
M7108 VDD 2763 2771 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=112370 $Y=16510 $D=111
M7109 2763 2762 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=112910 $Y=16510 $D=111
M7110 2765 2761 2763 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=113740 $Y=16260 $D=111
M7111 2774 2764 2765 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=114470 $Y=16260 $D=111
M7112 VDD 2767 2774 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=114800 $Y=16260 $D=111
M7113 2767 428 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=115260 $Y=16330 $D=111
M7114 VDD 2765 2767 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=115820 $Y=16040 $D=111
M7115 2766 2767 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=116430 $Y=16680 $D=111
M7116 VDD 2766 927 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=117370 $Y=16810 $D=111
M7117 result[13] 2767 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=117870 $Y=16810 $D=111
M7118 2785 287 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=109660 $Y=23480 $D=111
M7119 2778 2780 2785 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=109980 $Y=23480 $D=111
M7120 VDD 407 2778 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=110460 $Y=23480 $D=111
M7121 VDD clk 2777 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=110980 $Y=24070 $D=111
M7122 2780 2777 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=111490 $Y=24170 $D=111
M7123 2787 2777 2778 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=112050 $Y=23710 $D=111
M7124 VDD 2779 2787 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=112370 $Y=23710 $D=111
M7125 2779 2778 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=112910 $Y=23710 $D=111
M7126 2781 2777 2779 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=113740 $Y=23460 $D=111
M7127 2790 2780 2781 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=114470 $Y=23460 $D=111
M7128 VDD 2783 2790 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=114800 $Y=23460 $D=111
M7129 2783 407 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=115260 $Y=23530 $D=111
M7130 VDD 2781 2783 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=115820 $Y=23240 $D=111
M7131 2782 2783 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=116430 $Y=23880 $D=111
M7132 VDD 2782 928 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=117370 $Y=24010 $D=111
M7133 data_out[1] 2783 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=117870 $Y=24010 $D=111
M7134 2801 494 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=110060 $Y=50640 $D=111
M7135 2794 2796 2801 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=110380 $Y=50640 $D=111
M7136 VDD 425 2794 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=110860 $Y=50640 $D=111
M7137 VDD clk 2793 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=111380 $Y=49910 $D=111
M7138 2796 2793 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=111890 $Y=49950 $D=111
M7139 2803 2793 2794 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=112450 $Y=50410 $D=111
M7140 VDD 2795 2803 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=112770 $Y=50410 $D=111
M7141 2795 2794 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=113310 $Y=50410 $D=111
M7142 2797 2793 2795 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=114140 $Y=50660 $D=111
M7143 2806 2796 2797 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=114870 $Y=50660 $D=111
M7144 VDD 2799 2806 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=115200 $Y=50660 $D=111
M7145 2799 425 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=115660 $Y=50590 $D=111
M7146 VDD 2797 2799 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=116220 $Y=50880 $D=111
M7147 2798 2799 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=116830 $Y=50240 $D=111
M7148 VDD 2798 436 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=117770 $Y=50050 $D=111
M7149 839 2799 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=118270 $Y=50050 $D=111
M7150 2817 453 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=119260 $Y=21840 $D=111
M7151 2810 2812 2817 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=119580 $Y=21840 $D=111
M7152 VDD 428 2810 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=120060 $Y=21840 $D=111
M7153 VDD clk 2809 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=120580 $Y=21110 $D=111
M7154 2812 2809 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=121090 $Y=21150 $D=111
M7155 2819 2809 2810 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=121650 $Y=21610 $D=111
M7156 VDD 2811 2819 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=121970 $Y=21610 $D=111
M7157 2811 2810 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=122510 $Y=21610 $D=111
M7158 2813 2809 2811 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=123340 $Y=21860 $D=111
M7159 2822 2812 2813 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=124070 $Y=21860 $D=111
M7160 VDD 2815 2822 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=124400 $Y=21860 $D=111
M7161 2815 428 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=124860 $Y=21790 $D=111
M7162 VDD 2813 2815 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=125420 $Y=22080 $D=111
M7163 2814 2815 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=126030 $Y=21440 $D=111
M7164 VDD 2814 929 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=126970 $Y=21250 $D=111
M7165 result[14] 2815 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=127470 $Y=21250 $D=111
M7166 2833 398 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=132460 $Y=50640 $D=111
M7167 2826 2828 2833 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=132780 $Y=50640 $D=111
M7168 VDD 543 2826 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=133260 $Y=50640 $D=111
M7169 VDD clk 2825 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=133780 $Y=49910 $D=111
M7170 2828 2825 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=134290 $Y=49950 $D=111
M7171 2835 2825 2826 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=134850 $Y=50410 $D=111
M7172 VDD 2827 2835 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=135170 $Y=50410 $D=111
M7173 2827 2826 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=135710 $Y=50410 $D=111
M7174 2829 2825 2827 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=136540 $Y=50660 $D=111
M7175 2838 2828 2829 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=137270 $Y=50660 $D=111
M7176 VDD 2831 2838 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=137600 $Y=50660 $D=111
M7177 2831 543 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=138060 $Y=50590 $D=111
M7178 VDD 2829 2831 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=138620 $Y=50880 $D=111
M7179 2830 2831 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=139230 $Y=50240 $D=111
M7180 VDD 2830 930 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=140170 $Y=50050 $D=111
M7181 data_out[6] 2831 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=140670 $Y=50050 $D=111
M7182 2849 538 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=138460 $Y=52280 $D=111
M7183 2842 2844 2849 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=138780 $Y=52280 $D=111
M7184 VDD 544 2842 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=139260 $Y=52280 $D=111
M7185 VDD clk 2841 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=139780 $Y=52870 $D=111
M7186 2844 2841 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=140290 $Y=52970 $D=111
M7187 2851 2841 2842 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=140850 $Y=52510 $D=111
M7188 VDD 2843 2851 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=141170 $Y=52510 $D=111
M7189 2843 2842 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=141710 $Y=52510 $D=111
M7190 2845 2841 2843 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=142540 $Y=52260 $D=111
M7191 2854 2844 2845 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=143270 $Y=52260 $D=111
M7192 VDD 2847 2854 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=143600 $Y=52260 $D=111
M7193 2847 544 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=144060 $Y=52330 $D=111
M7194 VDD 2845 2847 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=144620 $Y=52040 $D=111
M7195 2846 2847 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=145230 $Y=52680 $D=111
M7196 VDD 2846 931 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=146170 $Y=52810 $D=111
M7197 data_out[7] 2847 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=146670 $Y=52810 $D=111
M7198 2865 367 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=141260 $Y=45080 $D=111
M7199 2858 2860 2865 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=141580 $Y=45080 $D=111
M7200 VDD 544 2858 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=142060 $Y=45080 $D=111
M7201 VDD clk 2857 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=142580 $Y=45670 $D=111
M7202 2860 2857 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=143090 $Y=45770 $D=111
M7203 2867 2857 2858 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=143650 $Y=45310 $D=111
M7204 VDD 2859 2867 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=143970 $Y=45310 $D=111
M7205 2859 2858 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=144510 $Y=45310 $D=111
M7206 2861 2857 2859 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=145340 $Y=45060 $D=111
M7207 2870 2860 2861 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=146070 $Y=45060 $D=111
M7208 VDD 2863 2870 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=146400 $Y=45060 $D=111
M7209 2863 544 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=146860 $Y=45130 $D=111
M7210 VDD 2861 2863 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=147420 $Y=44840 $D=111
M7211 2862 2863 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=148030 $Y=45480 $D=111
M7212 VDD 2862 932 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=148970 $Y=45610 $D=111
M7213 data_out[5] 2863 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=149470 $Y=45610 $D=111
M7214 2881 563 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=144060 $Y=21840 $D=111
M7215 2874 2876 2881 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=144380 $Y=21840 $D=111
M7216 VDD 564 2874 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=144860 $Y=21840 $D=111
M7217 VDD clk 2873 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=145380 $Y=21110 $D=111
M7218 2876 2873 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=145890 $Y=21150 $D=111
M7219 2883 2873 2874 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=146450 $Y=21610 $D=111
M7220 VDD 2875 2883 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=146770 $Y=21610 $D=111
M7221 2875 2874 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=147310 $Y=21610 $D=111
M7222 2877 2873 2875 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=148140 $Y=21860 $D=111
M7223 2886 2876 2877 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=148870 $Y=21860 $D=111
M7224 VDD 2879 2886 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=149200 $Y=21860 $D=111
M7225 2879 564 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=149660 $Y=21790 $D=111
M7226 VDD 2877 2879 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=150220 $Y=22080 $D=111
M7227 2878 2879 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=150830 $Y=21440 $D=111
M7228 VDD 2878 933 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=151770 $Y=21250 $D=111
M7229 result[24] 2879 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=152270 $Y=21250 $D=111
M7230 2897 176 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=144060 $Y=37880 $D=111
M7231 2890 2892 2897 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=144380 $Y=37880 $D=111
M7232 VDD 544 2890 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=144860 $Y=37880 $D=111
M7233 VDD clk 2889 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=145380 $Y=38470 $D=111
M7234 2892 2889 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=145890 $Y=38570 $D=111
M7235 2899 2889 2890 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=146450 $Y=38110 $D=111
M7236 VDD 2891 2899 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=146770 $Y=38110 $D=111
M7237 2891 2890 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=147310 $Y=38110 $D=111
M7238 2893 2889 2891 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=148140 $Y=37860 $D=111
M7239 2902 2892 2893 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=148870 $Y=37860 $D=111
M7240 VDD 2895 2902 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=149200 $Y=37860 $D=111
M7241 2895 544 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=149660 $Y=37930 $D=111
M7242 VDD 2893 2895 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=150220 $Y=37640 $D=111
M7243 2894 2895 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=150830 $Y=38280 $D=111
M7244 VDD 2894 934 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=151770 $Y=38410 $D=111
M7245 data_out[4] 2895 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=152270 $Y=38410 $D=111
M7246 2913 654 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=148060 $Y=23480 $D=111
M7247 2906 2908 2913 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=148380 $Y=23480 $D=111
M7248 VDD 662 2906 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=148860 $Y=23480 $D=111
M7249 VDD clk 2905 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=149380 $Y=24070 $D=111
M7250 2908 2905 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=149890 $Y=24170 $D=111
M7251 2915 2905 2906 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=150450 $Y=23710 $D=111
M7252 VDD 2907 2915 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=150770 $Y=23710 $D=111
M7253 2907 2906 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=151310 $Y=23710 $D=111
M7254 2909 2905 2907 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=152140 $Y=23460 $D=111
M7255 2918 2908 2909 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=152870 $Y=23460 $D=111
M7256 VDD 2911 2918 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=153200 $Y=23460 $D=111
M7257 2911 662 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=153660 $Y=23530 $D=111
M7258 VDD 2909 2911 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=154220 $Y=23240 $D=111
M7259 2910 2911 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=154830 $Y=23880 $D=111
M7260 VDD 2910 935 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=155770 $Y=24010 $D=111
M7261 result[23] 2911 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=156270 $Y=24010 $D=111
M7262 2929 621 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=156060 $Y=9080 $D=111
M7263 2922 2924 2929 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=156380 $Y=9080 $D=111
M7264 VDD 665 2922 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=156860 $Y=9080 $D=111
M7265 VDD clk 2921 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=157380 $Y=9670 $D=111
M7266 2924 2921 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=157890 $Y=9770 $D=111
M7267 2931 2921 2922 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=158450 $Y=9310 $D=111
M7268 VDD 2923 2931 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=158770 $Y=9310 $D=111
M7269 2923 2922 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=159310 $Y=9310 $D=111
M7270 2925 2921 2923 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=160140 $Y=9060 $D=111
M7271 2934 2924 2925 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=160870 $Y=9060 $D=111
M7272 VDD 2927 2934 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=161200 $Y=9060 $D=111
M7273 2927 665 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=161660 $Y=9130 $D=111
M7274 VDD 2925 2927 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=162220 $Y=8840 $D=111
M7275 2926 2927 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=162830 $Y=9480 $D=111
M7276 VDD 2926 936 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=163770 $Y=9610 $D=111
M7277 result[22] 2927 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=164270 $Y=9610 $D=111
M7278 2945 678 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=159660 $Y=21840 $D=111
M7279 2938 2940 2945 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=159980 $Y=21840 $D=111
M7280 VDD 638 2938 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=160460 $Y=21840 $D=111
M7281 VDD clk 2937 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=160980 $Y=21110 $D=111
M7282 2940 2937 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=161490 $Y=21150 $D=111
M7283 2947 2937 2938 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=162050 $Y=21610 $D=111
M7284 VDD 2939 2947 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=162370 $Y=21610 $D=111
M7285 2939 2938 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=162910 $Y=21610 $D=111
M7286 2941 2937 2939 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=163740 $Y=21860 $D=111
M7287 2950 2940 2941 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=164470 $Y=21860 $D=111
M7288 VDD 2943 2950 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=164800 $Y=21860 $D=111
M7289 2943 638 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=165260 $Y=21790 $D=111
M7290 VDD 2941 2943 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=165820 $Y=22080 $D=111
M7291 2942 2943 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=166430 $Y=21440 $D=111
M7292 VDD 2942 937 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=167370 $Y=21250 $D=111
M7293 result[27] 2943 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=167870 $Y=21250 $D=111
M7294 2961 643 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=160860 $Y=14640 $D=111
M7295 2954 2956 2961 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=161180 $Y=14640 $D=111
M7296 VDD 665 2954 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=161660 $Y=14640 $D=111
M7297 VDD clk 2953 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=162180 $Y=13910 $D=111
M7298 2956 2953 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=162690 $Y=13950 $D=111
M7299 2963 2953 2954 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=163250 $Y=14410 $D=111
M7300 VDD 2955 2963 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=163570 $Y=14410 $D=111
M7301 2955 2954 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=164110 $Y=14410 $D=111
M7302 2957 2953 2955 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=164940 $Y=14660 $D=111
M7303 2966 2956 2957 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=165670 $Y=14660 $D=111
M7304 VDD 2959 2966 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=166000 $Y=14660 $D=111
M7305 2959 665 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=166460 $Y=14590 $D=111
M7306 VDD 2957 2959 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=167020 $Y=14880 $D=111
M7307 2958 2959 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=167630 $Y=14240 $D=111
M7308 VDD 2958 938 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=168570 $Y=14050 $D=111
M7309 result[28] 2959 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=169070 $Y=14050 $D=111
M7310 2977 699 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=166460 $Y=9080 $D=111
M7311 2970 2972 2977 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=166780 $Y=9080 $D=111
M7312 VDD 665 2970 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=167260 $Y=9080 $D=111
M7313 VDD clk 2969 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=167780 $Y=9670 $D=111
M7314 2972 2969 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=168290 $Y=9770 $D=111
M7315 2979 2969 2970 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=168850 $Y=9310 $D=111
M7316 VDD 2971 2979 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=169170 $Y=9310 $D=111
M7317 2971 2970 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=169710 $Y=9310 $D=111
M7318 2973 2969 2971 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=170540 $Y=9060 $D=111
M7319 2982 2972 2973 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=171270 $Y=9060 $D=111
M7320 VDD 2975 2982 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=171600 $Y=9060 $D=111
M7321 2975 665 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=172060 $Y=9130 $D=111
M7322 VDD 2973 2975 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=172620 $Y=8840 $D=111
M7323 2974 2975 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=173230 $Y=9480 $D=111
M7324 VDD 2974 939 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=174170 $Y=9610 $D=111
M7325 result[29] 2975 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=174670 $Y=9610 $D=111
M7326 2993 708 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=168060 $Y=16280 $D=111
M7327 2986 2988 2993 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=168380 $Y=16280 $D=111
M7328 VDD 706 2986 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=168860 $Y=16280 $D=111
M7329 VDD clk 2985 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=169380 $Y=16870 $D=111
M7330 2988 2985 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=169890 $Y=16970 $D=111
M7331 2995 2985 2986 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=170450 $Y=16510 $D=111
M7332 VDD 2987 2995 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=170770 $Y=16510 $D=111
M7333 2987 2986 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=171310 $Y=16510 $D=111
M7334 2989 2985 2987 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=172140 $Y=16260 $D=111
M7335 2998 2988 2989 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=172870 $Y=16260 $D=111
M7336 VDD 2991 2998 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=173200 $Y=16260 $D=111
M7337 2991 706 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=173660 $Y=16330 $D=111
M7338 VDD 2989 2991 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=174220 $Y=16040 $D=111
M7339 2990 2991 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=174830 $Y=16680 $D=111
M7340 VDD 2990 940 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=175770 $Y=16810 $D=111
M7341 result[30] 2991 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=176270 $Y=16810 $D=111
M7342 3009 740 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=176060 $Y=9080 $D=111
M7343 3002 3004 3009 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=176380 $Y=9080 $D=111
M7344 VDD 665 3002 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=176860 $Y=9080 $D=111
M7345 VDD clk 3001 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=177380 $Y=9670 $D=111
M7346 3004 3001 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=177890 $Y=9770 $D=111
M7347 3011 3001 3002 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=178450 $Y=9310 $D=111
M7348 VDD 3003 3011 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=178770 $Y=9310 $D=111
M7349 3003 3002 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=179310 $Y=9310 $D=111
M7350 3005 3001 3003 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=180140 $Y=9060 $D=111
M7351 3014 3004 3005 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=180870 $Y=9060 $D=111
M7352 VDD 3007 3014 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=181200 $Y=9060 $D=111
M7353 3007 665 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=181660 $Y=9130 $D=111
M7354 VDD 3005 3007 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=182220 $Y=8840 $D=111
M7355 3006 3007 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=182830 $Y=9480 $D=111
M7356 VDD 3006 941 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=183770 $Y=9610 $D=111
M7357 result[31] 3007 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=184270 $Y=9610 $D=111
M7358 3018 80 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=18080 $Y=66790 $D=111
M7359 802 60 3018 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=18400 $Y=66790 $D=111
M7360 VDD 50 802 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=18920 $Y=66990 $D=111
M7361 3020 220 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=60480 $Y=57170 $D=111
M7362 229 215 3020 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=60800 $Y=57170 $D=111
M7363 VDD 210 229 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=61320 $Y=57170 $D=111
M7364 3022 412 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=110080 $Y=52390 $D=111
M7365 835 833 3022 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=110400 $Y=52390 $D=111
M7366 VDD 414 835 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=110920 $Y=52590 $D=111
M7367 3024 417 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=112080 $Y=64370 $D=111
M7368 420 435 3024 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=112400 $Y=64370 $D=111
M7369 VDD 476 420 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=112920 $Y=64370 $D=111
M7370 3026 458 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=121680 $Y=35570 $D=111
M7371 459 478 3026 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=122000 $Y=35570 $D=111
M7372 VDD 477 459 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=122520 $Y=35570 $D=111
M7373 3028 492 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=131280 $Y=37990 $D=111
M7374 506 502 3028 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=131600 $Y=37990 $D=111
M7375 VDD 517 506 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=132120 $Y=38190 $D=111
M7376 3030 522 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=135280 $Y=30790 $D=111
M7377 546 527 3030 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=135600 $Y=30790 $D=111
M7378 VDD 551 546 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=136120 $Y=30990 $D=111
M7379 3032 528 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=137280 $Y=30790 $D=111
M7380 537 530 3032 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=137600 $Y=30790 $D=111
M7381 VDD 536 537 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=138120 $Y=30990 $D=111
M7382 3034 600 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=146080 $Y=49970 $D=111
M7383 606 587 3034 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=146400 $Y=49970 $D=111
M7384 VDD 580 606 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=146920 $Y=49970 $D=111
M7385 3036 581 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=146480 $Y=57170 $D=111
M7386 559 566 3036 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=146800 $Y=57170 $D=111
M7387 VDD 607 559 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=147320 $Y=57170 $D=111
M7388 3038 591 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=147280 $Y=35570 $D=111
M7389 596 571 3038 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=147600 $Y=35570 $D=111
M7390 VDD 585 596 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=148120 $Y=35570 $D=111
M7391 3040 626 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=156080 $Y=59590 $D=111
M7392 687 616 3040 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=156400 $Y=59590 $D=111
M7393 VDD 627 687 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=156920 $Y=59790 $D=111
M7394 3042 783 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=174880 $Y=59590 $D=111
M7395 775 784 3042 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=175200 $Y=59590 $D=111
M7396 VDD 736 775 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=175720 $Y=59790 $D=111
M7397 3044 703 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=4.172e-13 pd=1.04e-06 ps=3.18e-06 nrd=0.119048 nrs=0.59127 sa=3.7e-07 sb=1.06667e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=175680 $Y=49970 $D=111
M7398 727 721 3044 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.81622e-13 as=8.4e-14 pd=1.40757e-06 ps=1.04e-06 nrd=0.2574 nrs=0.119048 sa=6.9e-07 sb=7.46667e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=176000 $Y=49970 $D=111
M7399 VDD 724 727 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.984e-13 as=1.38378e-13 pd=3.2e-06 ps=1.07243e-06 nrd=0.972656 nrs=0.337838 sa=1.21e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=176520 $Y=49970 $D=111
M7400 22 70 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=4.47266e-13 pd=3.24e-06 ps=3.17595e-06 nrd=0.246154 nrs=0.264654 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=17830 $Y=30390 $D=111
M7401 204 167 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=4.47266e-13 pd=3.24e-06 ps=3.17595e-06 nrd=0.246154 nrs=0.264654 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=51030 $Y=15990 $D=111
M7402 286 285 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=4.47266e-13 pd=3.24e-06 ps=3.17595e-06 nrd=0.246154 nrs=0.264654 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=75830 $Y=42710 $D=111
M7403 830 353 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=4.47266e-13 pd=3.24e-06 ps=3.17595e-06 nrd=0.246154 nrs=0.264654 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=95430 $Y=71510 $D=111
M7404 584 850 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=4.47266e-13 pd=3.24e-06 ps=3.17595e-06 nrd=0.246154 nrs=0.264654 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=139830 $Y=13910 $D=111
M7405 719 674 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=4.47266e-13 pd=3.24e-06 ps=3.17595e-06 nrd=0.246154 nrs=0.264654 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=175430 $Y=71510 $D=111
M7406 112 89 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.42e-13 pd=1.66e-06 ps=3.28e-06 nrd=0.138462 nrs=0.261538 sa=3.4e-07 sb=1.31662e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=27300 $Y=42710 $D=111
M7407 VDD 89 112 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.39919e-13 as=2.34e-13 pd=1.75447e-06 ps=1.66e-06 nrd=0.141964 nrs=0.138462 sa=8.2e-07 sb=8.36615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=27780 $Y=42710 $D=111
M7408 112 89 VDD VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.944e-13 as=2.14081e-13 pd=3.18e-06 ps=1.56553e-06 nrd=0.36742 nrs=0.159097 sa=1.3e-06 sb=4.26207e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=28260 $Y=42710 $D=111
M7409 201 172 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.42e-13 pd=1.66e-06 ps=3.28e-06 nrd=0.138462 nrs=0.261538 sa=3.4e-07 sb=1.31662e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=50900 $Y=73590 $D=111
M7410 VDD 172 201 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.39919e-13 as=2.34e-13 pd=1.75447e-06 ps=1.66e-06 nrd=0.141964 nrs=0.138462 sa=8.2e-07 sb=8.36615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=51380 $Y=73590 $D=111
M7411 201 172 VDD VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.944e-13 as=2.14081e-13 pd=3.18e-06 ps=1.56553e-06 nrd=0.36742 nrs=0.159097 sa=1.3e-06 sb=4.26207e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=51860 $Y=73730 $D=111
M7412 263 201 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.42e-13 pd=1.66e-06 ps=3.28e-06 nrd=0.138462 nrs=0.261538 sa=3.4e-07 sb=1.31662e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=60900 $Y=49910 $D=111
M7413 VDD 201 263 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.39919e-13 as=2.34e-13 pd=1.75447e-06 ps=1.66e-06 nrd=0.141964 nrs=0.138462 sa=8.2e-07 sb=8.36615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=61380 $Y=49910 $D=111
M7414 263 201 VDD VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.944e-13 as=2.14081e-13 pd=3.18e-06 ps=1.56553e-06 nrd=0.36742 nrs=0.159097 sa=1.3e-06 sb=4.26207e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=61860 $Y=49910 $D=111
M7415 518 849 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.42e-13 pd=1.66e-06 ps=3.28e-06 nrd=0.138462 nrs=0.261538 sa=3.4e-07 sb=1.31662e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=134100 $Y=64310 $D=111
M7416 VDD 849 518 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.39919e-13 as=2.34e-13 pd=1.75447e-06 ps=1.66e-06 nrd=0.141964 nrs=0.138462 sa=8.2e-07 sb=8.36615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=134580 $Y=64310 $D=111
M7417 518 849 VDD VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.944e-13 as=2.14081e-13 pd=3.18e-06 ps=1.56553e-06 nrd=0.36742 nrs=0.159097 sa=1.3e-06 sb=4.26207e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=135060 $Y=64310 $D=111
M7418 562 849 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.42e-13 pd=1.66e-06 ps=3.28e-06 nrd=0.138462 nrs=0.261538 sa=3.4e-07 sb=1.31662e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=135300 $Y=66390 $D=111
M7419 VDD 849 562 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.39919e-13 as=2.34e-13 pd=1.75447e-06 ps=1.66e-06 nrd=0.141964 nrs=0.138462 sa=8.2e-07 sb=8.36615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=135780 $Y=66390 $D=111
M7420 562 849 VDD VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.944e-13 as=2.14081e-13 pd=3.18e-06 ps=1.56553e-06 nrd=0.36742 nrs=0.159097 sa=1.3e-06 sb=4.26207e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=136260 $Y=66530 $D=111
M7421 742 523 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.42e-13 pd=1.66e-06 ps=3.28e-06 nrd=0.138462 nrs=0.261538 sa=3.4e-07 sb=1.31662e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=169300 $Y=35510 $D=111
M7422 VDD 523 742 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.39919e-13 as=2.34e-13 pd=1.75447e-06 ps=1.66e-06 nrd=0.141964 nrs=0.138462 sa=8.2e-07 sb=8.36615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=169780 $Y=35510 $D=111
M7423 742 523 VDD VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.944e-13 as=2.14081e-13 pd=3.18e-06 ps=1.56553e-06 nrd=0.36742 nrs=0.159097 sa=1.3e-06 sb=4.26207e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=170260 $Y=35510 $D=111
M7424 729 523 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.42e-13 pd=1.66e-06 ps=3.28e-06 nrd=0.138462 nrs=0.261538 sa=3.4e-07 sb=1.31662e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=173300 $Y=64310 $D=111
M7425 VDD 523 729 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.39919e-13 as=2.34e-13 pd=1.75447e-06 ps=1.66e-06 nrd=0.141964 nrs=0.138462 sa=8.2e-07 sb=8.36615e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=173780 $Y=64310 $D=111
M7426 729 523 VDD VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.944e-13 as=2.14081e-13 pd=3.18e-06 ps=1.56553e-06 nrd=0.36742 nrs=0.159097 sa=1.3e-06 sb=4.26207e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=174260 $Y=64310 $D=111
M7427 3046 85 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.90476e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=25920 $Y=71510 $D=111
M7428 885 81 3046 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.82857e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=26240 $Y=71510 $D=111
M7429 3047 81 885 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=1.59238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=26720 $Y=71510 $D=111
M7430 VDD 85 3047 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.57903e-13 as=8.4e-14 pd=1.58919e-06 ps=1.04e-06 nrd=0.365508 nrs=0.119048 sa=1.44e-06 sb=1.27238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=27040 $Y=71510 $D=111
M7431 885 91 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.96497e-13 pd=1e-06 ps=1.21081e-06 nrd=0.28125 nrs=0.47973 sa=2e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=27720 $Y=71510 $D=111
M7432 VDD 91 885 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.41426e-13 as=1.152e-13 pd=2.68522e-06 ps=1e-06 nrd=0.83356 nrs=0.28125 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=28200 $Y=71510 $D=111
M7433 3049 218 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.90476e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=58320 $Y=52450 $D=111
M7434 220 221 3049 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.82857e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=58640 $Y=52450 $D=111
M7435 3050 221 220 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=1.59238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=59120 $Y=52450 $D=111
M7436 VDD 218 3050 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.57903e-13 as=8.4e-14 pd=1.58919e-06 ps=1.04e-06 nrd=0.365508 nrs=0.119048 sa=1.44e-06 sb=1.27238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=59440 $Y=52450 $D=111
M7437 220 247 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.96497e-13 pd=1e-06 ps=1.21081e-06 nrd=0.28125 nrs=0.47973 sa=2e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=60120 $Y=52650 $D=111
M7438 VDD 247 220 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.41426e-13 as=1.152e-13 pd=2.68522e-06 ps=1e-06 nrd=0.83356 nrs=0.28125 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=60600 $Y=52650 $D=111
M7439 3052 281 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.90476e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=63120 $Y=21110 $D=111
M7440 235 249 3052 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.82857e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=63440 $Y=21110 $D=111
M7441 3053 249 235 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=1.59238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=63920 $Y=21110 $D=111
M7442 VDD 281 3053 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.57903e-13 as=8.4e-14 pd=1.58919e-06 ps=1.04e-06 nrd=0.365508 nrs=0.119048 sa=1.44e-06 sb=1.27238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=64240 $Y=21110 $D=111
M7443 235 258 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.96497e-13 pd=1e-06 ps=1.21081e-06 nrd=0.28125 nrs=0.47973 sa=2e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=64920 $Y=21110 $D=111
M7444 VDD 258 235 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.41426e-13 as=1.152e-13 pd=2.68522e-06 ps=1e-06 nrd=0.83356 nrs=0.28125 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=65400 $Y=21110 $D=111
M7445 3055 439 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.90476e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=116720 $Y=71510 $D=111
M7446 840 435 3055 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.82857e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=117040 $Y=71510 $D=111
M7447 3056 435 840 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=1.59238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=117520 $Y=71510 $D=111
M7448 VDD 439 3056 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.57903e-13 as=8.4e-14 pd=1.58919e-06 ps=1.04e-06 nrd=0.365508 nrs=0.119048 sa=1.44e-06 sb=1.27238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=117840 $Y=71510 $D=111
M7449 840 468 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.96497e-13 pd=1e-06 ps=1.21081e-06 nrd=0.28125 nrs=0.47973 sa=2e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=118520 $Y=71510 $D=111
M7450 VDD 468 840 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.41426e-13 as=1.152e-13 pd=2.68522e-06 ps=1e-06 nrd=0.83356 nrs=0.28125 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=119000 $Y=71510 $D=111
M7451 3058 574 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.90476e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=157520 $Y=57110 $D=111
M7452 664 637 3058 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.82857e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=157840 $Y=57110 $D=111
M7453 3059 637 664 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=1.59238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=158320 $Y=57110 $D=111
M7454 VDD 574 3059 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.57903e-13 as=8.4e-14 pd=1.58919e-06 ps=1.04e-06 nrd=0.365508 nrs=0.119048 sa=1.44e-06 sb=1.27238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=158640 $Y=57110 $D=111
M7455 664 649 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.96497e-13 pd=1e-06 ps=1.21081e-06 nrd=0.28125 nrs=0.47973 sa=2e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=159320 $Y=57110 $D=111
M7456 VDD 649 664 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.41426e-13 as=1.152e-13 pd=2.68522e-06 ps=1e-06 nrd=0.83356 nrs=0.28125 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=159800 $Y=57110 $D=111
M7457 3061 648 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.90476e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=158720 $Y=59650 $D=111
M7458 674 659 3061 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.82857e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=159040 $Y=59650 $D=111
M7459 3062 659 674 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=1.59238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=159520 $Y=59650 $D=111
M7460 VDD 648 3062 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.57903e-13 as=8.4e-14 pd=1.58919e-06 ps=1.04e-06 nrd=0.365508 nrs=0.119048 sa=1.44e-06 sb=1.27238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=159840 $Y=59650 $D=111
M7461 674 640 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.96497e-13 pd=1e-06 ps=1.21081e-06 nrd=0.28125 nrs=0.47973 sa=2e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=160520 $Y=59850 $D=111
M7462 VDD 640 674 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.41426e-13 as=1.152e-13 pd=2.68522e-06 ps=1e-06 nrd=0.83356 nrs=0.28125 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=161000 $Y=59850 $D=111
M7463 3064 686 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.90476e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=171120 $Y=66850 $D=111
M7464 758 719 3064 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.82857e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=171440 $Y=66850 $D=111
M7465 3065 719 758 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=1.59238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=171920 $Y=66850 $D=111
M7466 VDD 686 3065 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.57903e-13 as=8.4e-14 pd=1.58919e-06 ps=1.04e-06 nrd=0.365508 nrs=0.119048 sa=1.44e-06 sb=1.27238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=172240 $Y=66850 $D=111
M7467 758 692 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.96497e-13 pd=1e-06 ps=1.21081e-06 nrd=0.28125 nrs=0.47973 sa=2e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=172920 $Y=67050 $D=111
M7468 VDD 692 758 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.41426e-13 as=1.152e-13 pd=2.68522e-06 ps=1e-06 nrd=0.83356 nrs=0.28125 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=173400 $Y=67050 $D=111
M7469 3067 731 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=1.90476e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=173120 $Y=38050 $D=111
M7470 741 690 3067 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=1.82857e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=173440 $Y=38050 $D=111
M7471 3068 690 741 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.12e-06 sb=1.59238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=173920 $Y=38050 $D=111
M7472 VDD 731 3068 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.57903e-13 as=8.4e-14 pd=1.58919e-06 ps=1.04e-06 nrd=0.365508 nrs=0.119048 sa=1.44e-06 sb=1.27238e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=174240 $Y=38050 $D=111
M7473 741 735 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.96497e-13 pd=1e-06 ps=1.21081e-06 nrd=0.28125 nrs=0.47973 sa=2e-06 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=174920 $Y=38250 $D=111
M7474 VDD 735 741 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.41426e-13 as=1.152e-13 pd=2.68522e-06 ps=1e-06 nrd=0.83356 nrs=0.28125 sa=2e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=175400 $Y=38250 $D=111
M7475 3069 69 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.06e-13 as=3.392e-13 pd=1.26e-06 ps=2.76e-06 nrd=0.0943396 nrs=0.301887 sa=3.2e-07 sb=1.84151e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=22210 $Y=64310 $D=111
M7476 80 121 3069 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04512e-13 as=1.06e-13 pd=1.55596e-06 ps=1.26e-06 nrd=0.182015 nrs=0.0943396 sa=6.4e-07 sb=1.73434e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=22530 $Y=64310 $D=111
M7477 3070 121 80 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.16088e-13 pd=1.32e-06 ps=1.64404e-06 nrd=0.0892857 nrs=0.172264 sa=9.83393e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=23010 $Y=64430 $D=111
M7478 VDD 69 3070 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.30339e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=23330 $Y=64430 $D=111
M7479 3071 69 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.78339e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=23810 $Y=64430 $D=111
M7480 80 121 3071 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=1.90196e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=24130 $Y=64430 $D=111
M7481 3072 125 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.06e-13 as=3.392e-13 pd=1.26e-06 ps=2.76e-06 nrd=0.0943396 nrs=0.301887 sa=3.2e-07 sb=1.84151e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=35410 $Y=28310 $D=111
M7482 119 130 3072 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04512e-13 as=1.06e-13 pd=1.55596e-06 ps=1.26e-06 nrd=0.182015 nrs=0.0943396 sa=6.4e-07 sb=1.73434e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=35730 $Y=28310 $D=111
M7483 3073 130 119 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.16088e-13 pd=1.32e-06 ps=1.64404e-06 nrd=0.0892857 nrs=0.172264 sa=9.83393e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=36210 $Y=28430 $D=111
M7484 VDD 125 3073 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.30339e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=36530 $Y=28430 $D=111
M7485 3074 125 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.78339e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=37010 $Y=28430 $D=111
M7486 119 130 3074 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=1.90196e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=37330 $Y=28430 $D=111
M7487 3075 191 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.06e-13 as=3.392e-13 pd=1.26e-06 ps=2.76e-06 nrd=0.0943396 nrs=0.301887 sa=3.2e-07 sb=1.84151e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=37010 $Y=73830 $D=111
M7488 81 238 3075 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04512e-13 as=1.06e-13 pd=1.55596e-06 ps=1.26e-06 nrd=0.182015 nrs=0.0943396 sa=6.4e-07 sb=1.73434e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=37330 $Y=73830 $D=111
M7489 3076 238 81 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.16088e-13 pd=1.32e-06 ps=1.64404e-06 nrd=0.0892857 nrs=0.172264 sa=9.83393e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=37810 $Y=73650 $D=111
M7490 VDD 191 3076 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.30339e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=38130 $Y=73650 $D=111
M7491 3077 191 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.78339e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=38610 $Y=73650 $D=111
M7492 81 238 3077 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=1.90196e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=38930 $Y=73650 $D=111
M7493 3078 308 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.06e-13 as=3.392e-13 pd=1.26e-06 ps=2.76e-06 nrd=0.0943396 nrs=0.301887 sa=3.2e-07 sb=1.84151e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=82210 $Y=73830 $D=111
M7494 366 347 3078 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04512e-13 as=1.06e-13 pd=1.55596e-06 ps=1.26e-06 nrd=0.182015 nrs=0.0943396 sa=6.4e-07 sb=1.73434e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=82530 $Y=73830 $D=111
M7495 3079 347 366 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.16088e-13 pd=1.32e-06 ps=1.64404e-06 nrd=0.0892857 nrs=0.172264 sa=9.83393e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=83010 $Y=73650 $D=111
M7496 VDD 308 3079 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.30339e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=83330 $Y=73650 $D=111
M7497 3080 308 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.78339e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=83810 $Y=73650 $D=111
M7498 366 347 3080 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=1.90196e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=84130 $Y=73650 $D=111
M7499 3081 353 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.06e-13 as=3.392e-13 pd=1.26e-06 ps=2.76e-06 nrd=0.0943396 nrs=0.301887 sa=3.2e-07 sb=1.84151e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=92610 $Y=73830 $D=111
M7500 473 366 3081 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04512e-13 as=1.06e-13 pd=1.55596e-06 ps=1.26e-06 nrd=0.182015 nrs=0.0943396 sa=6.4e-07 sb=1.73434e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=92930 $Y=73830 $D=111
M7501 3082 366 473 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.16088e-13 pd=1.32e-06 ps=1.64404e-06 nrd=0.0892857 nrs=0.172264 sa=9.83393e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=93410 $Y=73650 $D=111
M7502 VDD 353 3082 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.30339e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=93730 $Y=73650 $D=111
M7503 3083 353 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.78339e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=94210 $Y=73650 $D=111
M7504 473 366 3083 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=1.90196e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=94530 $Y=73650 $D=111
M7505 3084 846 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.06e-13 as=3.392e-13 pd=1.26e-06 ps=2.76e-06 nrd=0.0943396 nrs=0.301887 sa=3.2e-07 sb=1.84151e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=127010 $Y=71510 $D=111
M7506 490 417 3084 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04512e-13 as=1.06e-13 pd=1.55596e-06 ps=1.26e-06 nrd=0.182015 nrs=0.0943396 sa=6.4e-07 sb=1.73434e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=127330 $Y=71510 $D=111
M7507 3085 417 490 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.16088e-13 pd=1.32e-06 ps=1.64404e-06 nrd=0.0892857 nrs=0.172264 sa=9.83393e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=127810 $Y=71630 $D=111
M7508 VDD 846 3085 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.30339e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=128130 $Y=71630 $D=111
M7509 3086 846 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.78339e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=128610 $Y=71630 $D=111
M7510 490 417 3086 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=1.90196e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=128930 $Y=71630 $D=111
M7511 3087 485 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.06e-13 as=3.392e-13 pd=1.26e-06 ps=2.76e-06 nrd=0.0943396 nrs=0.301887 sa=3.2e-07 sb=1.84151e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=130210 $Y=57110 $D=111
M7512 508 521 3087 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04512e-13 as=1.06e-13 pd=1.55596e-06 ps=1.26e-06 nrd=0.182015 nrs=0.0943396 sa=6.4e-07 sb=1.73434e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=130530 $Y=57110 $D=111
M7513 3088 521 508 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.16088e-13 pd=1.32e-06 ps=1.64404e-06 nrd=0.0892857 nrs=0.172264 sa=9.83393e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=131010 $Y=57230 $D=111
M7514 VDD 485 3088 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.30339e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=131330 $Y=57230 $D=111
M7515 3089 485 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.78339e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=131810 $Y=57230 $D=111
M7516 508 521 3089 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=1.90196e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=132130 $Y=57230 $D=111
M7517 3090 681 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.06e-13 as=3.392e-13 pd=1.26e-06 ps=2.76e-06 nrd=0.0943396 nrs=0.301887 sa=3.2e-07 sb=1.84151e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=168610 $Y=42710 $D=111
M7518 694 700 3090 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04512e-13 as=1.06e-13 pd=1.55596e-06 ps=1.26e-06 nrd=0.182015 nrs=0.0943396 sa=6.4e-07 sb=1.73434e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=168930 $Y=42710 $D=111
M7519 3091 700 694 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.16088e-13 pd=1.32e-06 ps=1.64404e-06 nrd=0.0892857 nrs=0.172264 sa=9.83393e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=169410 $Y=42830 $D=111
M7520 VDD 681 3091 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.30339e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=169730 $Y=42830 $D=111
M7521 3092 681 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.78339e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=170210 $Y=42830 $D=111
M7522 694 700 3092 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=1.90196e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=170530 $Y=42830 $D=111
M7523 3093 693 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.06e-13 as=3.392e-13 pd=1.26e-06 ps=2.76e-06 nrd=0.0943396 nrs=0.301887 sa=3.2e-07 sb=1.84151e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=172210 $Y=23430 $D=111
M7524 704 743 3093 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04512e-13 as=1.06e-13 pd=1.55596e-06 ps=1.26e-06 nrd=0.182015 nrs=0.0943396 sa=6.4e-07 sb=1.73434e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=172530 $Y=23430 $D=111
M7525 3094 743 704 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.16088e-13 pd=1.32e-06 ps=1.64404e-06 nrd=0.0892857 nrs=0.172264 sa=9.83393e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=173010 $Y=23250 $D=111
M7526 VDD 693 3094 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.30339e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=173330 $Y=23250 $D=111
M7527 3095 693 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.78339e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=173810 $Y=23250 $D=111
M7528 704 743 3095 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=1.90196e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=174130 $Y=23250 $D=111
M7529 3096 581 VDD VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.4e-14 as=1.408e-13 pd=6.4e-07 ps=1.52e-06 nrd=0.227273 nrs=0.727273 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=142160 $Y=60050 $D=111
M7530 556 557 3096 VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=4.4e-14 pd=1.52e-06 ps=6.4e-07 nrd=0.727273 nrs=0.227273 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=142480 $Y=60050 $D=111
M7531 3097 666 VDD VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.4e-14 as=1.408e-13 pd=6.4e-07 ps=1.52e-06 nrd=0.227273 nrs=0.727273 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=164160 $Y=57110 $D=111
M7532 653 667 3097 VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=4.4e-14 pd=1.52e-06 ps=6.4e-07 nrd=0.727273 nrs=0.227273 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=164480 $Y=57110 $D=111
M7533 3098 713 VDD VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.4e-14 as=1.408e-13 pd=6.4e-07 ps=1.52e-06 nrd=0.227273 nrs=0.727273 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=165760 $Y=57110 $D=111
M7534 691 667 3098 VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=4.4e-14 pd=1.52e-06 ps=6.4e-07 nrd=0.727273 nrs=0.227273 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=166080 $Y=57110 $D=111
M7535 3099 683 VDD VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.4e-14 as=1.408e-13 pd=6.4e-07 ps=1.52e-06 nrd=0.227273 nrs=0.727273 sa=3.2e-07 sb=6.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=171760 $Y=35510 $D=111
M7536 731 709 3099 VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.408e-13 as=4.4e-14 pd=1.52e-06 ps=6.4e-07 nrd=0.727273 nrs=0.227273 sa=6.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=172080 $Y=35510 $D=111
M7537 VDD 14 3100 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=15210 $Y=52440 $D=111
M7538 3100 13 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=15690 $Y=52440 $D=111
M7539 45 38 3100 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=16170 $Y=52440 $D=111
M7540 VDD 443 3102 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=123610 $Y=66840 $D=111
M7541 3102 465 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=124090 $Y=66840 $D=111
M7542 468 467 3102 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=124570 $Y=66840 $D=111
M7543 VDD 484 3104 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=128810 $Y=30840 $D=111
M7544 3104 501 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=129290 $Y=30840 $D=111
M7545 527 847 3104 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=129770 $Y=30840 $D=111
M7546 VDD 515 3106 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=128810 $Y=35520 $D=111
M7547 3106 506 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=129290 $Y=35520 $D=111
M7548 530 851 3106 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=129770 $Y=35520 $D=111
M7549 VDD 914 3108 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=140410 $Y=30840 $D=111
M7550 3108 558 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=140890 $Y=30840 $D=111
M7551 551 550 3108 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=141370 $Y=30840 $D=111
M7552 VDD 601 3110 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=150410 $Y=52440 $D=111
M7553 3110 598 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=150890 $Y=52440 $D=111
M7554 566 619 3110 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=151370 $Y=52440 $D=111
M7555 VDD 599 3112 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=151210 $Y=59640 $D=111
M7556 3112 602 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=151690 $Y=59640 $D=111
M7557 627 603 3112 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=152170 $Y=59640 $D=111
M7558 VDD 635 3114 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=154010 $Y=57120 $D=111
M7559 3114 625 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=154490 $Y=57120 $D=111
M7560 616 629 3114 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=154970 $Y=57120 $D=111
M7561 VDD 685 3116 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=168810 $Y=57120 $D=111
M7562 3116 687 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=169290 $Y=57120 $D=111
M7563 721 718 3116 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=169770 $Y=57120 $D=111
M7564 VDD 862 3118 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=170810 $Y=57120 $D=111
M7565 3118 684 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=171290 $Y=57120 $D=111
M7566 725 698 3118 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=171770 $Y=57120 $D=111
M7567 VDD 773 3120 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=2.688e-13 pd=1.2e-06 ps=2.32e-06 nrd=0.214286 nrs=0.380952 sa=3.2e-07 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=171210 $Y=59640 $D=111
M7568 3120 732 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=1.512e-13 pd=1.2e-06 ps=1.2e-06 nrd=0.214286 nrs=0.214286 sa=8e-07 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=171690 $Y=59640 $D=111
M7569 714 747 3120 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.688e-13 as=1.512e-13 pd=2.32e-06 ps=1.2e-06 nrd=0.380952 nrs=0.214286 sa=1.28e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=172170 $Y=59640 $D=111
M7570 VDD weight_in[1] 3122 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85906e-13 as=3.264e-13 pd=1.45461e-06 ps=2.68e-06 nrd=0.178687 nrs=0.313725 sa=3.2e-07 sb=1.32e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=25800 $Y=73850 $D=111
M7571 86 3122 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.33294e-13 pd=1.64e-06 ps=1.82539e-06 nrd=0.140625 nrs=0.142391 sa=6.78125e-07 sb=8.4e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=26280 $Y=73590 $D=111
M7572 VDD 3122 86 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.40123e-13 as=2.304e-13 pd=3.13436e-06 ps=1.64e-06 nrd=0.26863 nrs=0.140625 sa=1.15813e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=26760 $Y=73590 $D=111
M7573 VDD 101 3123 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85906e-13 as=3.264e-13 pd=1.45461e-06 ps=2.68e-06 nrd=0.178687 nrs=0.313725 sa=3.2e-07 sb=1.32e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=29400 $Y=28330 $D=111
M7574 129 3123 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.33294e-13 pd=1.64e-06 ps=1.82539e-06 nrd=0.140625 nrs=0.142391 sa=6.78125e-07 sb=8.4e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=29880 $Y=28330 $D=111
M7575 VDD 3123 129 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.40123e-13 as=2.304e-13 pd=3.13436e-06 ps=1.64e-06 nrd=0.26863 nrs=0.140625 sa=1.15813e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=30360 $Y=28330 $D=111
M7576 VDD 127 3124 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85906e-13 as=3.264e-13 pd=1.45461e-06 ps=2.68e-06 nrd=0.178687 nrs=0.313725 sa=3.2e-07 sb=1.32e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=31000 $Y=35530 $D=111
M7577 192 3124 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.33294e-13 pd=1.64e-06 ps=1.82539e-06 nrd=0.140625 nrs=0.142391 sa=6.78125e-07 sb=8.4e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=31480 $Y=35530 $D=111
M7578 VDD 3124 192 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.40123e-13 as=2.304e-13 pd=3.13436e-06 ps=1.64e-06 nrd=0.26863 nrs=0.140625 sa=1.15813e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=31960 $Y=35530 $D=111
M7579 VDD 98 3125 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85906e-13 as=3.264e-13 pd=1.45461e-06 ps=2.68e-06 nrd=0.178687 nrs=0.313725 sa=3.2e-07 sb=1.32e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=37800 $Y=59450 $D=111
M7580 151 3125 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.33294e-13 pd=1.64e-06 ps=1.82539e-06 nrd=0.140625 nrs=0.142391 sa=6.78125e-07 sb=8.4e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=38280 $Y=59190 $D=111
M7581 VDD 3125 151 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.40123e-13 as=2.304e-13 pd=3.13436e-06 ps=1.64e-06 nrd=0.26863 nrs=0.140625 sa=1.15813e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=38760 $Y=59190 $D=111
M7582 VDD 187 3126 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85906e-13 as=3.264e-13 pd=1.45461e-06 ps=2.68e-06 nrd=0.178687 nrs=0.313725 sa=3.2e-07 sb=1.32e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=69800 $Y=45050 $D=111
M7583 283 3126 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.33294e-13 pd=1.64e-06 ps=1.82539e-06 nrd=0.140625 nrs=0.142391 sa=6.78125e-07 sb=8.4e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=70280 $Y=44790 $D=111
M7584 VDD 3126 283 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.40123e-13 as=2.304e-13 pd=3.13436e-06 ps=1.64e-06 nrd=0.26863 nrs=0.140625 sa=1.15813e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=70760 $Y=44790 $D=111
M7585 VDD 263 3127 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85906e-13 as=3.264e-13 pd=1.45461e-06 ps=2.68e-06 nrd=0.178687 nrs=0.313725 sa=3.2e-07 sb=1.32e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=70600 $Y=35530 $D=111
M7586 170 3127 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.33294e-13 pd=1.64e-06 ps=1.82539e-06 nrd=0.140625 nrs=0.142391 sa=6.78125e-07 sb=8.4e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=71080 $Y=35530 $D=111
M7587 VDD 3127 170 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.40123e-13 as=2.304e-13 pd=3.13436e-06 ps=1.64e-06 nrd=0.26863 nrs=0.140625 sa=1.15813e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=71560 $Y=35530 $D=111
M7588 VDD 263 3128 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85906e-13 as=3.264e-13 pd=1.45461e-06 ps=2.68e-06 nrd=0.178687 nrs=0.313725 sa=3.2e-07 sb=1.32e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=72600 $Y=45050 $D=111
M7589 307 3128 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.33294e-13 pd=1.64e-06 ps=1.82539e-06 nrd=0.140625 nrs=0.142391 sa=6.78125e-07 sb=8.4e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=73080 $Y=44790 $D=111
M7590 VDD 3128 307 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.40123e-13 as=2.304e-13 pd=3.13436e-06 ps=1.64e-06 nrd=0.26863 nrs=0.140625 sa=1.15813e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=73560 $Y=44790 $D=111
M7591 VDD 171 3129 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85906e-13 as=3.264e-13 pd=1.45461e-06 ps=2.68e-06 nrd=0.178687 nrs=0.313725 sa=3.2e-07 sb=1.32e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=102600 $Y=49930 $D=111
M7592 398 3129 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.33294e-13 pd=1.64e-06 ps=1.82539e-06 nrd=0.140625 nrs=0.142391 sa=6.78125e-07 sb=8.4e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=103080 $Y=49930 $D=111
M7593 VDD 3129 398 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.40123e-13 as=2.304e-13 pd=3.13436e-06 ps=1.64e-06 nrd=0.26863 nrs=0.140625 sa=1.15813e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=103560 $Y=49930 $D=111
M7594 VDD 584 3130 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85906e-13 as=3.264e-13 pd=1.45461e-06 ps=2.68e-06 nrd=0.178687 nrs=0.313725 sa=3.2e-07 sb=1.32e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=148200 $Y=16250 $D=111
M7595 638 3130 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.33294e-13 pd=1.64e-06 ps=1.82539e-06 nrd=0.140625 nrs=0.142391 sa=6.78125e-07 sb=8.4e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=148680 $Y=15990 $D=111
M7596 VDD 3130 638 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.40123e-13 as=2.304e-13 pd=3.13436e-06 ps=1.64e-06 nrd=0.26863 nrs=0.140625 sa=1.15813e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=149160 $Y=15990 $D=111
M7597 VDD 641 3131 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.85906e-13 as=3.264e-13 pd=1.45461e-06 ps=2.68e-06 nrd=0.178687 nrs=0.313725 sa=3.2e-07 sb=1.32e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=170600 $Y=30650 $D=111
M7598 706 3131 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.33294e-13 pd=1.64e-06 ps=1.82539e-06 nrd=0.140625 nrs=0.142391 sa=6.78125e-07 sb=8.4e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=171080 $Y=30390 $D=111
M7599 VDD 3131 706 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.40123e-13 as=2.304e-13 pd=3.13436e-06 ps=1.64e-06 nrd=0.26863 nrs=0.140625 sa=1.15813e-06 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=171560 $Y=30390 $D=111
M7600 VDD 11 3132 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-14 panw9=2.16e-14 panw10=0 $X=8980 $Y=31150 $D=111
M7601 23 3132 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-13 $X=9470 $Y=30390 $D=111
M7602 VDD data_in[4] 3133 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-14 panw9=2.16e-14 panw10=0 $X=8980 $Y=49910 $D=111
M7603 136 3133 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-13 $X=9470 $Y=49910 $D=111
M7604 VDD data_in[6] 3134 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-14 panw9=2.16e-14 panw10=0 $X=8980 $Y=59950 $D=111
M7605 797 3134 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-13 $X=9470 $Y=59190 $D=111
M7606 VDD data_in[3] 3135 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=10980 $Y=35510 $D=111
M7607 127 3135 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=11470 $Y=35510 $D=111
M7608 VDD 85 3136 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=13380 $Y=67150 $D=111
M7609 50 3136 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=13870 $Y=66390 $D=111
M7610 VDD rst_n 3137 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=19380 $Y=74350 $D=111
M7611 32 3137 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=19870 $Y=73590 $D=111
M7612 VDD 803 3138 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=23380 $Y=71510 $D=111
M7613 58 3138 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=23870 $Y=71510 $D=111
M7614 VDD 131 3139 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=46580 $Y=49910 $D=111
M7615 180 3139 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=47070 $Y=49910 $D=111
M7616 VDD 128 3140 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=5.4e-14 $X=48580 $Y=9550 $D=111
M7617 202 3140 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.52e-14 panw8=4.8e-14 panw9=9.6e-14 panw10=9.6e-14 $X=49070 $Y=8790 $D=111
M7618 VDD 129 3141 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=58580 $Y=23950 $D=111
M7619 217 3141 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=59070 $Y=23190 $D=111
M7620 VDD 271 3142 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=61380 $Y=21110 $D=111
M7621 11 3142 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=61870 $Y=21110 $D=111
M7622 VDD 187 3143 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=63380 $Y=49910 $D=111
M7623 241 3143 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=63870 $Y=49910 $D=111
M7624 VDD 202 3144 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=64980 $Y=13910 $D=111
M7625 252 3144 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=65470 $Y=13910 $D=111
M7626 VDD 256 3145 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=71780 $Y=21110 $D=111
M7627 271 3145 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=72270 $Y=21110 $D=111
M7628 VDD 49 3146 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=73780 $Y=23950 $D=111
M7629 287 3146 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=74270 $Y=23190 $D=111
M7630 VDD 318 3147 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=82580 $Y=21110 $D=111
M7631 256 3147 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=83070 $Y=21110 $D=111
M7632 VDD 303 3148 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=85780 $Y=31150 $D=111
M7633 329 3148 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=86270 $Y=30390 $D=111
M7634 VDD 186 3149 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=86980 $Y=52750 $D=111
M7635 538 3149 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=87470 $Y=51990 $D=111
M7636 VDD 358 3150 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=97780 $Y=64310 $D=111
M7637 376 3150 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=98270 $Y=64310 $D=111
M7638 VDD 399 3151 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=105380 $Y=16750 $D=111
M7639 389 3151 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=105870 $Y=15990 $D=111
M7640 VDD 407 3152 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=106580 $Y=31150 $D=111
M7641 425 3152 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=107070 $Y=30390 $D=111
M7642 VDD 407 3153 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=108180 $Y=23950 $D=111
M7643 374 3153 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=108670 $Y=23190 $D=111
M7644 VDD 409 3154 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=108580 $Y=52750 $D=111
M7645 437 3154 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=109070 $Y=51990 $D=111
M7646 VDD 437 3155 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=117780 $Y=57110 $D=111
M7647 485 3155 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=118270 $Y=57110 $D=111
M7648 VDD 396 3156 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=121780 $Y=16750 $D=111
M7649 526 3156 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=122270 $Y=15990 $D=111
M7650 VDD 425 3157 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=124980 $Y=57110 $D=111
M7651 543 3157 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=125470 $Y=57110 $D=111
M7652 VDD 526 3158 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=135380 $Y=13910 $D=111
M7653 570 3158 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=135870 $Y=13910 $D=111
M7654 VDD 500 3159 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=141780 $Y=16750 $D=111
M7655 611 3159 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=142270 $Y=15990 $D=111
M7656 VDD 611 3160 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=147780 $Y=28310 $D=111
M7657 582 3160 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=148270 $Y=28310 $D=111
M7658 VDD 697 3161 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=152580 $Y=52750 $D=111
M7659 610 3161 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=153070 $Y=51990 $D=111
M7660 VDD 611 3162 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=153380 $Y=16750 $D=111
M7661 593 3162 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=153870 $Y=15990 $D=111
M7662 VDD 638 3163 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=159380 $Y=13910 $D=111
M7663 665 3163 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=159870 $Y=13910 $D=111
M7664 VDD 645 3164 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=161780 $Y=16750 $D=111
M7665 701 3164 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=162270 $Y=15990 $D=111
M7666 VDD 682 3165 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=169380 $Y=23950 $D=111
M7667 688 3165 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=169870 $Y=23190 $D=111
M7668 VDD data_in[1] 3166 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=5.52e-14 panw8=8.64e-14 panw9=9.6e-15 panw10=0 $X=8820 $Y=28310 $D=111
M7669 49 3166 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.08e-13 panw10=3.84e-14 $X=9380 $Y=28310 $D=111
M7670 VDD 3166 49 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=1.152e-13 $X=9860 $Y=28310 $D=111
M7671 VDD 797 3167 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=5.52e-14 panw8=8.64e-14 panw9=9.6e-15 panw10=0 $X=8820 $Y=57110 $D=111
M7672 171 3167 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.08e-13 panw10=3.84e-14 $X=9380 $Y=57110 $D=111
M7673 VDD 3167 171 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=1.152e-13 $X=9860 $Y=57110 $D=111
M7674 VDD 32 3168 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=20020 $Y=57110 $D=111
M7675 68 3168 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=20580 $Y=57110 $D=111
M7676 VDD 3168 68 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=21060 $Y=57110 $D=111
M7677 VDD weight_in[0] 3169 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=22420 $Y=74110 $D=111
M7678 97 3169 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=22980 $Y=73930 $D=111
M7679 VDD 3169 97 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=23460 $Y=73930 $D=111
M7680 VDD 82 3170 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=23620 $Y=35510 $D=111
M7681 74 3170 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=24180 $Y=35510 $D=111
M7682 VDD 3170 74 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=24660 $Y=35510 $D=111
M7683 VDD weight_in[2] 3171 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=28020 $Y=74110 $D=111
M7684 79 3171 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=28580 $Y=73930 $D=111
M7685 VDD 3171 79 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=29060 $Y=73930 $D=111
M7686 VDD 73 3172 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=30420 $Y=59710 $D=111
M7687 189 3172 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=30980 $Y=59530 $D=111
M7688 VDD 3172 189 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=31460 $Y=59530 $D=111
M7689 VDD 211 3173 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=36820 $Y=64310 $D=111
M7690 139 3173 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=37380 $Y=64310 $D=111
M7691 VDD 3173 139 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=37860 $Y=64310 $D=111
M7692 VDD weight_in[4] 3174 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=36820 $Y=71510 $D=111
M7693 153 3174 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=37380 $Y=71510 $D=111
M7694 VDD 3174 153 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=37860 $Y=71510 $D=111
M7695 VDD weight_in[5] 3175 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=44420 $Y=74110 $D=111
M7696 172 3175 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=44980 $Y=73930 $D=111
M7697 VDD 3175 172 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=45460 $Y=73930 $D=111
M7698 VDD weight_in[7] 3176 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=48820 $Y=74110 $D=111
M7699 187 3176 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=49380 $Y=73930 $D=111
M7700 VDD 3176 187 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=49860 $Y=73930 $D=111
M7701 VDD 141 3177 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=53620 $Y=30910 $D=111
M7702 254 3177 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=54180 $Y=30730 $D=111
M7703 VDD 3177 254 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=54660 $Y=30730 $D=111
M7704 VDD 213 3178 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=56020 $Y=52510 $D=111
M7705 218 3178 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=56580 $Y=52330 $D=111
M7706 VDD 3178 218 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=57060 $Y=52330 $D=111
M7707 VDD fire_in 3179 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=57620 $Y=74110 $D=111
M7708 306 3179 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=58180 $Y=73930 $D=111
M7709 VDD 3179 306 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=58660 $Y=73930 $D=111
M7710 VDD 187 3180 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=65220 $Y=42710 $D=111
M7711 240 3180 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=65780 $Y=42710 $D=111
M7712 VDD 3180 240 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=66260 $Y=42710 $D=111
M7713 VDD 252 3181 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=68020 $Y=13910 $D=111
M7714 299 3181 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=68580 $Y=13910 $D=111
M7715 VDD 3181 299 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=69060 $Y=13910 $D=111
M7716 VDD 246 3182 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=78420 $Y=57110 $D=111
M7717 295 3182 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=78980 $Y=57110 $D=111
M7718 VDD 3182 295 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=79460 $Y=57110 $D=111
M7719 VDD 157 3183 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=93620 $Y=38110 $D=111
M7720 367 3183 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=94180 $Y=37930 $D=111
M7721 VDD 3183 367 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=94660 $Y=37930 $D=111
M7722 VDD 348 3184 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=94820 $Y=57110 $D=111
M7723 360 3184 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=95380 $Y=57110 $D=111
M7724 VDD 3184 360 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=95860 $Y=57110 $D=111
M7725 VDD 371 3185 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=7.2e-14 $X=114820 $Y=9310 $D=111
M7726 428 3185 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6.36e-14 panw10=7.2e-14 $X=115380 $Y=9130 $D=111
M7727 VDD 3185 428 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=6.36e-14 panw10=7.2e-14 $X=115860 $Y=9130 $D=111
M7728 VDD 408 3186 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=123220 $Y=16510 $D=111
M7729 491 3186 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=123780 $Y=16330 $D=111
M7730 VDD 3186 491 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=124260 $Y=16330 $D=111
M7731 VDD 428 3187 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=125220 $Y=16510 $D=111
M7732 479 3187 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=125780 $Y=16330 $D=111
M7733 VDD 3187 479 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=126260 $Y=16330 $D=111
M7734 VDD 491 3188 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=129220 $Y=13910 $D=111
M7735 500 3188 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=129780 $Y=13910 $D=111
M7736 VDD 3188 500 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=130260 $Y=13910 $D=111
M7737 VDD 638 3189 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=164420 $Y=23710 $D=111
M7738 662 3189 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=164980 $Y=23530 $D=111
M7739 VDD 3189 662 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=165460 $Y=23530 $D=111
M7740 VDD 689 3190 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82897e-13 as=2.496e-13 pd=1.25517e-06 ps=2.2e-06 nrd=0.300619 nrs=0.410256 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=167620 $Y=28310 $D=111
M7741 693 3190 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=2.25103e-13 pd=1.32e-06 ps=1.54483e-06 nrd=0.1875 nrs=0.244253 sa=7.825e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=168180 $Y=28310 $D=111
M7742 VDD 3190 693 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.168e-13 as=1.728e-13 pd=2.58e-06 ps=1.32e-06 nrd=0.34375 nrs=0.1875 sa=1.2625e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=168660 $Y=28310 $D=111
M7743 27 26 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=16120 $Y=28310 $D=111
M7744 47 62 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=17320 $Y=28310 $D=111
M7745 76 117 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=23320 $Y=13910 $D=111
M7746 117 68 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=24520 $Y=13910 $D=111
M7747 303 302 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=78920 $Y=21110 $D=111
M7748 302 299 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=80120 $Y=21110 $D=111
M7749 344 316 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=93720 $Y=13910 $D=111
M7750 356 344 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=94920 $Y=13910 $D=111
M7751 525 492 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=134520 $Y=42710 $D=111
M7752 912 517 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=135720 $Y=42710 $D=111
M7753 534 502 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=136920 $Y=57110 $D=111
M7754 586 485 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=138120 $Y=57110 $D=111
M7755 655 620 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=157320 $Y=21110 $D=111
M7756 645 655 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=158520 $Y=21110 $D=111
M7757 658 662 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=159320 $Y=30410 $D=111
M7758 641 658 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=160520 $Y=30410 $D=111
M7759 667 669 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=163320 $Y=49910 $D=111
M7760 659 598 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=164520 $Y=49910 $D=111
M7761 860 688 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=166920 $Y=30410 $D=111
M7762 681 860 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.44718e-13 pd=3.2e-06 ps=3.16718e-06 nrd=0.25 nrs=0.271434 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=168120 $Y=30410 $D=111
M7763 VDD clk 3191 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02606e-13 as=1.792e-13 pd=1.02366e-06 ps=1.76e-06 nrd=0.327189 nrs=0.571429 sa=3.2e-07 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=119280 $Y=49910 $D=111
M7764 3199 clk VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.83219e-13 as=2.38194e-13 pd=1.60469e-06 ps=2.37634e-06 nrd=0.108413 nrs=0.140943 sa=4.51692e-07 sb=6.15385e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=119680 $Y=49910 $D=111
M7765 3195 3196 3199 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.88e-13 as=1.77581e-13 pd=3.16e-06 ps=1.55531e-06 nrd=0.181406 nrs=0.111855 sa=8.55873e-07 sb=2.28571e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=120080 $Y=49910 $D=111
M7766 VDD 508 3192 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41429e-13 as=2.112e-13 pd=1.18446e-06 ps=1.96e-06 nrd=0.324675 nrs=0.484848 sa=3.2e-07 sb=1.38667e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=120900 $Y=49910 $D=111
M7767 3196 3191 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.40816e-13 as=2.78571e-13 pd=2.09515e-06 ps=2.33304e-06 nrd=0.142494 nrs=0.164835 sa=5.34462e-07 sb=1.13046e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=121340 $Y=49910 $D=111
M7768 VDD 3191 3196 VDD lppfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46635e-13 as=1.40784e-13 pd=1.36353e-06 ps=1.22485e-06 nrd=0.25387 nrs=0.24374 sa=1.02263e-06 sb=1.64842e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=121820 $Y=50130 $D=111
M7769 3200 3196 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.85224e-13 pd=1.16e-06 ps=1.72235e-06 nrd=0.104167 nrs=0.20098 sa=1.02958e-06 sb=1.48e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=122260 $Y=50250 $D=111
M7770 3193 3192 3200 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=9.6e-14 pd=1.32e-06 ps=1.16e-06 nrd=0.1875 nrs=0.104167 sa=1.34958e-06 sb=1.16e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=122580 $Y=50250 $D=111
M7771 3202 3192 3193 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.728e-13 pd=1.16e-06 ps=1.32e-06 nrd=0.104167 nrs=0.1875 sa=1.66875e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=123060 $Y=50250 $D=111
M7772 VDD 3196 3202 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.2609e-13 as=9.6e-14 pd=2.46194e-06 ps=1.16e-06 nrd=0.353831 nrs=0.104167 sa=1.78833e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=123380 $Y=50250 $D=111
M7773 3204 3195 3193 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.008e-13 pd=4.8e-07 ps=1.28e-06 nrd=0.357143 nrs=1.28571 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1e-15 panw8=1.6e-14 panw9=1.66e-14 panw10=0 $X=124580 $Y=50490 $D=111
M7774 VDD 3194 3204 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.95304e-14 as=2.8e-14 pd=6.05652e-07 ps=4.8e-07 nrd=0.759317 nrs=0.357143 sa=6.8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.44e-14 panw9=1.92e-14 panw10=0 $X=124900 $Y=50490 $D=111
M7775 3194 3193 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.72139e-13 pd=1.64e-06 ps=2.7687e-06 nrd=0.140625 nrs=0.166101 sa=4.21562e-07 sb=1.42e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=125340 $Y=49930 $D=111
M7776 VDD 3193 3194 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.48524e-13 as=2.304e-13 pd=2.25416e-06 ps=1.64e-06 nrd=0.151687 nrs=0.140625 sa=9.01562e-07 sb=1.2025e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=125820 $Y=49930 $D=111
M7777 3194 543 VDD VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.35912e-13 pd=1.06e-06 ps=1.23274e-06 nrd=0.257143 nrs=0.27737 sa=1.47429e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=126260 $Y=50110 $D=111
M7778 3198 3195 3194 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.76229e-06 sb=1.73771e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=126740 $Y=50110 $D=111
M7779 3194 3195 3198 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=1.25771e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=127220 $Y=50110 $D=111
M7780 3198 3195 3194 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=7.77714e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=127700 $Y=50110 $D=111
M7781 3194 3195 3198 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.084e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.425306 nrs=0.257143 sa=2e-06 sb=2.97714e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=128180 $Y=50110 $D=111
M7782 3210 3197 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.779e-13 pd=4.8e-07 ps=2.32e-06 nrd=0.357143 nrs=3.54464 sa=4.3e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.2e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=129310 $Y=50510 $D=111
M7783 3198 3196 3210 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.24e-14 as=2.8e-14 pd=6.34286e-07 ps=4.8e-07 nrd=0.923469 nrs=0.357143 sa=7.5e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=5e-15 panw8=1.6e-14 panw9=1.26e-14 panw10=0 $X=129630 $Y=50510 $D=111
M7784 VDD 543 3198 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.72667e-13 as=1.81e-13 pd=1.21579e-06 ps=1.58571e-06 nrd=0.352381 nrs=0.369388 sa=7.1e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.2e-14 panw9=4.8e-14 panw10=2.4e-14 $X=130160 $Y=50510 $D=111
M7785 VDD 3198 3197 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.90667e-14 as=1.064e-13 pd=4.86316e-07 ps=1.32e-06 nrd=0.880952 nrs=1.35714 sa=3.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=130480 $Y=49910 $D=111
M7786 456 3198 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=3.20667e-13 pd=1.66e-06 ps=2.25789e-06 nrd=0.138462 nrs=0.189744 sa=9.87231e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=130880 $Y=49910 $D=111
M7787 VDD 3198 456 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.34e-13 pd=3.24e-06 ps=1.66e-06 nrd=0.246154 nrs=0.138462 sa=1.36385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=131360 $Y=49910 $D=111
M7788 VDD clk 3211 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02606e-13 as=1.792e-13 pd=1.02366e-06 ps=1.76e-06 nrd=0.327189 nrs=0.571429 sa=3.2e-07 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=140480 $Y=42710 $D=111
M7789 3219 clk VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.83219e-13 as=2.38194e-13 pd=1.60469e-06 ps=2.37634e-06 nrd=0.108413 nrs=0.140943 sa=4.51692e-07 sb=6.15385e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=140880 $Y=42710 $D=111
M7790 3215 3216 3219 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.88e-13 as=1.77581e-13 pd=3.16e-06 ps=1.55531e-06 nrd=0.181406 nrs=0.111855 sa=8.55873e-07 sb=2.28571e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=141280 $Y=42710 $D=111
M7791 VDD 540 3212 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41429e-13 as=2.112e-13 pd=1.18446e-06 ps=1.96e-06 nrd=0.324675 nrs=0.484848 sa=3.2e-07 sb=1.38667e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=142100 $Y=42710 $D=111
M7792 3216 3211 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.40816e-13 as=2.78571e-13 pd=2.09515e-06 ps=2.33304e-06 nrd=0.142494 nrs=0.164835 sa=5.34462e-07 sb=1.13046e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=142540 $Y=42710 $D=111
M7793 VDD 3211 3216 VDD lppfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46635e-13 as=1.40784e-13 pd=1.36353e-06 ps=1.22485e-06 nrd=0.25387 nrs=0.24374 sa=1.02263e-06 sb=1.64842e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=143020 $Y=42930 $D=111
M7794 3220 3216 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.85224e-13 pd=1.16e-06 ps=1.72235e-06 nrd=0.104167 nrs=0.20098 sa=1.02958e-06 sb=1.48e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=143460 $Y=43050 $D=111
M7795 3213 3212 3220 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=9.6e-14 pd=1.32e-06 ps=1.16e-06 nrd=0.1875 nrs=0.104167 sa=1.34958e-06 sb=1.16e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=143780 $Y=43050 $D=111
M7796 3222 3212 3213 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.728e-13 pd=1.16e-06 ps=1.32e-06 nrd=0.104167 nrs=0.1875 sa=1.66875e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=144260 $Y=43050 $D=111
M7797 VDD 3216 3222 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.2609e-13 as=9.6e-14 pd=2.46194e-06 ps=1.16e-06 nrd=0.353831 nrs=0.104167 sa=1.78833e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=144580 $Y=43050 $D=111
M7798 3224 3215 3213 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.008e-13 pd=4.8e-07 ps=1.28e-06 nrd=0.357143 nrs=1.28571 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1e-15 panw8=1.6e-14 panw9=1.66e-14 panw10=0 $X=145780 $Y=43290 $D=111
M7799 VDD 3214 3224 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.95304e-14 as=2.8e-14 pd=6.05652e-07 ps=4.8e-07 nrd=0.759317 nrs=0.357143 sa=6.8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.44e-14 panw9=1.92e-14 panw10=0 $X=146100 $Y=43290 $D=111
M7800 3214 3213 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.72139e-13 pd=1.64e-06 ps=2.7687e-06 nrd=0.140625 nrs=0.166101 sa=4.21562e-07 sb=1.42e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=146540 $Y=42730 $D=111
M7801 VDD 3213 3214 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.48524e-13 as=2.304e-13 pd=2.25416e-06 ps=1.64e-06 nrd=0.151687 nrs=0.140625 sa=9.01562e-07 sb=1.2025e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=147020 $Y=42730 $D=111
M7802 3214 564 VDD VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.35912e-13 pd=1.06e-06 ps=1.23274e-06 nrd=0.257143 nrs=0.27737 sa=1.47429e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=147460 $Y=42910 $D=111
M7803 3218 3215 3214 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.76229e-06 sb=1.73771e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=147940 $Y=42910 $D=111
M7804 3214 3215 3218 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=1.25771e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=148420 $Y=42910 $D=111
M7805 3218 3215 3214 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=7.77714e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=148900 $Y=42910 $D=111
M7806 3214 3215 3218 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.084e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.425306 nrs=0.257143 sa=2e-06 sb=2.97714e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=149380 $Y=42910 $D=111
M7807 3230 3217 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.779e-13 pd=4.8e-07 ps=2.32e-06 nrd=0.357143 nrs=3.54464 sa=4.3e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.2e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=150510 $Y=43310 $D=111
M7808 3218 3216 3230 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.24e-14 as=2.8e-14 pd=6.34286e-07 ps=4.8e-07 nrd=0.923469 nrs=0.357143 sa=7.5e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=5e-15 panw8=1.6e-14 panw9=1.26e-14 panw10=0 $X=150830 $Y=43310 $D=111
M7809 VDD 564 3218 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.72667e-13 as=1.81e-13 pd=1.21579e-06 ps=1.58571e-06 nrd=0.352381 nrs=0.369388 sa=7.1e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.2e-14 panw9=4.8e-14 panw10=2.4e-14 $X=151360 $Y=43310 $D=111
M7810 VDD 3218 3217 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.90667e-14 as=1.064e-13 pd=4.86316e-07 ps=1.32e-06 nrd=0.880952 nrs=1.35714 sa=3.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=151680 $Y=42710 $D=111
M7811 568 3218 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=3.20667e-13 pd=1.66e-06 ps=2.25789e-06 nrd=0.138462 nrs=0.189744 sa=9.87231e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=152080 $Y=42710 $D=111
M7812 VDD 3218 568 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.34e-13 pd=3.24e-06 ps=1.66e-06 nrd=0.246154 nrs=0.138462 sa=1.36385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=152560 $Y=42710 $D=111
M7813 VDD clk 3231 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02606e-13 as=1.792e-13 pd=1.02366e-06 ps=1.76e-06 nrd=0.327189 nrs=0.571429 sa=3.2e-07 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=146880 $Y=74330 $D=111
M7814 3239 clk VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.83219e-13 as=2.38194e-13 pd=1.60469e-06 ps=2.37634e-06 nrd=0.108413 nrs=0.140943 sa=4.51692e-07 sb=6.15385e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=147280 $Y=73590 $D=111
M7815 3235 3236 3239 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.88e-13 as=1.77581e-13 pd=3.16e-06 ps=1.55531e-06 nrd=0.181406 nrs=0.111855 sa=8.55873e-07 sb=2.28571e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=147680 $Y=73630 $D=111
M7816 VDD 856 3232 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41429e-13 as=2.112e-13 pd=1.18446e-06 ps=1.96e-06 nrd=0.324675 nrs=0.484848 sa=3.2e-07 sb=1.38667e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=148500 $Y=74230 $D=111
M7817 3236 3231 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.40816e-13 as=2.78571e-13 pd=2.09515e-06 ps=2.33304e-06 nrd=0.142494 nrs=0.164835 sa=5.34462e-07 sb=1.13046e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=148940 $Y=73590 $D=111
M7818 VDD 3231 3236 VDD lppfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46635e-13 as=1.40784e-13 pd=1.36353e-06 ps=1.22485e-06 nrd=0.25387 nrs=0.24374 sa=1.02263e-06 sb=1.64842e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=149420 $Y=73910 $D=111
M7819 3240 3236 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.85224e-13 pd=1.16e-06 ps=1.72235e-06 nrd=0.104167 nrs=0.20098 sa=1.02958e-06 sb=1.48e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=149860 $Y=73590 $D=111
M7820 3233 3232 3240 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=9.6e-14 pd=1.32e-06 ps=1.16e-06 nrd=0.1875 nrs=0.104167 sa=1.34958e-06 sb=1.16e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=150180 $Y=73590 $D=111
M7821 3242 3232 3233 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.728e-13 pd=1.16e-06 ps=1.32e-06 nrd=0.104167 nrs=0.1875 sa=1.66875e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=150660 $Y=73590 $D=111
M7822 VDD 3236 3242 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.2609e-13 as=9.6e-14 pd=2.46194e-06 ps=1.16e-06 nrd=0.353831 nrs=0.104167 sa=1.78833e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=150980 $Y=73590 $D=111
M7823 3244 3235 3233 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.008e-13 pd=4.8e-07 ps=1.28e-06 nrd=0.357143 nrs=1.28571 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1e-15 panw8=1.6e-14 panw9=1.66e-14 panw10=0 $X=152180 $Y=74030 $D=111
M7824 VDD 3234 3244 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.95304e-14 as=2.8e-14 pd=6.05652e-07 ps=4.8e-07 nrd=0.759317 nrs=0.357143 sa=6.8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.44e-14 panw9=1.92e-14 panw10=0 $X=152500 $Y=74030 $D=111
M7825 3234 3233 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.72139e-13 pd=1.64e-06 ps=2.7687e-06 nrd=0.140625 nrs=0.166101 sa=4.21562e-07 sb=1.42e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=152940 $Y=73590 $D=111
M7826 VDD 3233 3234 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.48524e-13 as=2.304e-13 pd=2.25416e-06 ps=1.64e-06 nrd=0.151687 nrs=0.140625 sa=9.01562e-07 sb=1.2025e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=153420 $Y=73590 $D=111
M7827 3234 610 VDD VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.35912e-13 pd=1.06e-06 ps=1.23274e-06 nrd=0.257143 nrs=0.27737 sa=1.47429e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=153860 $Y=73990 $D=111
M7828 3238 3235 3234 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.76229e-06 sb=1.73771e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=154340 $Y=73990 $D=111
M7829 3234 3235 3238 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=1.25771e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=154820 $Y=73990 $D=111
M7830 3238 3235 3234 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=7.77714e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=155300 $Y=73990 $D=111
M7831 3234 3235 3238 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.084e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.425306 nrs=0.257143 sa=2e-06 sb=2.97714e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=155780 $Y=73990 $D=111
M7832 3250 3237 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.779e-13 pd=4.8e-07 ps=2.32e-06 nrd=0.357143 nrs=3.54464 sa=4.3e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.2e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=156910 $Y=74010 $D=111
M7833 3238 3236 3250 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.24e-14 as=2.8e-14 pd=6.34286e-07 ps=4.8e-07 nrd=0.923469 nrs=0.357143 sa=7.5e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=5e-15 panw8=1.6e-14 panw9=1.26e-14 panw10=0 $X=157230 $Y=74010 $D=111
M7834 VDD 610 3238 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.72667e-13 as=1.81e-13 pd=1.21579e-06 ps=1.58571e-06 nrd=0.352381 nrs=0.369388 sa=7.1e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.2e-14 panw9=4.8e-14 panw10=2.4e-14 $X=157760 $Y=73590 $D=111
M7835 VDD 3238 3237 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.90667e-14 as=1.064e-13 pd=4.86316e-07 ps=1.32e-06 nrd=0.880952 nrs=1.35714 sa=3.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=158080 $Y=74610 $D=111
M7836 609 3238 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=3.20667e-13 pd=1.66e-06 ps=2.25789e-06 nrd=0.138462 nrs=0.189744 sa=9.87231e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=158480 $Y=73590 $D=111
M7837 VDD 3238 609 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.34e-13 pd=3.24e-06 ps=1.66e-06 nrd=0.246154 nrs=0.138462 sa=1.36385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=158960 $Y=73590 $D=111
M7838 VDD clk 3251 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.02606e-13 as=1.792e-13 pd=1.02366e-06 ps=1.76e-06 nrd=0.327189 nrs=0.571429 sa=3.2e-07 sb=1e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=164880 $Y=52730 $D=111
M7839 3259 clk VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.83219e-13 as=2.38194e-13 pd=1.60469e-06 ps=2.37634e-06 nrd=0.108413 nrs=0.140943 sa=4.51692e-07 sb=6.15385e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=165280 $Y=51990 $D=111
M7840 3255 3256 3259 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.88e-13 as=1.77581e-13 pd=3.16e-06 ps=1.55531e-06 nrd=0.181406 nrs=0.111855 sa=8.55873e-07 sb=2.28571e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=165680 $Y=52030 $D=111
M7841 VDD 664 3252 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.41429e-13 as=2.112e-13 pd=1.18446e-06 ps=1.96e-06 nrd=0.324675 nrs=0.484848 sa=3.2e-07 sb=1.38667e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=166500 $Y=52630 $D=111
M7842 3256 3251 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.40816e-13 as=2.78571e-13 pd=2.09515e-06 ps=2.33304e-06 nrd=0.142494 nrs=0.164835 sa=5.34462e-07 sb=1.13046e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=166940 $Y=51990 $D=111
M7843 VDD 3251 3256 VDD lppfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.46635e-13 as=1.40784e-13 pd=1.36353e-06 ps=1.22485e-06 nrd=0.25387 nrs=0.24374 sa=1.02263e-06 sb=1.64842e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=167420 $Y=52310 $D=111
M7844 3260 3256 VDD VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.85224e-13 pd=1.16e-06 ps=1.72235e-06 nrd=0.104167 nrs=0.20098 sa=1.02958e-06 sb=1.48e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=167860 $Y=51990 $D=111
M7845 3253 3252 3260 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.728e-13 as=9.6e-14 pd=1.32e-06 ps=1.16e-06 nrd=0.1875 nrs=0.104167 sa=1.34958e-06 sb=1.16e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=168180 $Y=51990 $D=111
M7846 3262 3252 3253 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.728e-13 pd=1.16e-06 ps=1.32e-06 nrd=0.104167 nrs=0.1875 sa=1.66875e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=168660 $Y=51990 $D=111
M7847 VDD 3256 3262 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.2609e-13 as=9.6e-14 pd=2.46194e-06 ps=1.16e-06 nrd=0.353831 nrs=0.104167 sa=1.78833e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=8.4e-15 $X=168980 $Y=51990 $D=111
M7848 3264 3255 3253 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.008e-13 pd=4.8e-07 ps=1.28e-06 nrd=0.357143 nrs=1.28571 sa=3.6e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1e-15 panw8=1.6e-14 panw9=1.66e-14 panw10=0 $X=170180 $Y=52430 $D=111
M7849 VDD 3254 3264 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.95304e-14 as=2.8e-14 pd=6.05652e-07 ps=4.8e-07 nrd=0.759317 nrs=0.357143 sa=6.8e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.44e-14 panw9=1.92e-14 panw10=0 $X=170500 $Y=52430 $D=111
M7850 3254 3253 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.72139e-13 pd=1.64e-06 ps=2.7687e-06 nrd=0.140625 nrs=0.166101 sa=4.21562e-07 sb=1.42e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=170940 $Y=51990 $D=111
M7851 VDD 3253 3254 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.48524e-13 as=2.304e-13 pd=2.25416e-06 ps=1.64e-06 nrd=0.151687 nrs=0.140625 sa=9.01562e-07 sb=1.2025e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=171420 $Y=51990 $D=111
M7852 3254 697 VDD VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.35912e-13 pd=1.06e-06 ps=1.23274e-06 nrd=0.257143 nrs=0.27737 sa=1.47429e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=171860 $Y=52390 $D=111
M7853 3258 3255 3254 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=1.76229e-06 sb=1.73771e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=172340 $Y=52390 $D=111
M7854 3254 3255 3258 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=1.25771e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=172820 $Y=52390 $D=111
M7855 3258 3255 3254 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26e-13 as=1.26e-13 pd=1.06e-06 ps=1.06e-06 nrd=0.257143 nrs=0.257143 sa=2e-06 sb=7.77714e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=173300 $Y=52390 $D=111
M7856 3254 3255 3258 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.084e-13 as=1.26e-13 pd=2.04e-06 ps=1.06e-06 nrd=0.425306 nrs=0.257143 sa=2e-06 sb=2.97714e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=173780 $Y=52390 $D=111
M7857 3270 3257 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.779e-13 pd=4.8e-07 ps=2.32e-06 nrd=0.357143 nrs=3.54464 sa=4.3e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.2e-14 panw8=2.16e-14 panw9=0 panw10=0 $X=174910 $Y=52410 $D=111
M7858 3258 3256 3270 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.24e-14 as=2.8e-14 pd=6.34286e-07 ps=4.8e-07 nrd=0.923469 nrs=0.357143 sa=7.5e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=5e-15 panw8=1.6e-14 panw9=1.26e-14 panw10=0 $X=175230 $Y=52410 $D=111
M7859 VDD 697 3258 VDD lppfet w=7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.72667e-13 as=1.81e-13 pd=1.21579e-06 ps=1.58571e-06 nrd=0.352381 nrs=0.369388 sa=7.1e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.2e-14 panw9=4.8e-14 panw10=2.4e-14 $X=175760 $Y=51990 $D=111
M7860 VDD 3258 3257 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.90667e-14 as=1.064e-13 pd=4.86316e-07 ps=1.32e-06 nrd=0.880952 nrs=1.35714 sa=3.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=176080 $Y=53010 $D=111
M7861 597 3258 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=3.20667e-13 pd=1.66e-06 ps=2.25789e-06 nrd=0.138462 nrs=0.189744 sa=9.87231e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=176480 $Y=51990 $D=111
M7862 VDD 3258 597 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.34e-13 pd=3.24e-06 ps=1.66e-06 nrd=0.246154 nrs=0.138462 sa=1.36385e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=176960 $Y=51990 $D=111
M7863 VDD data_in[5] 3271 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-14 panw9=2.16e-14 panw10=0 $X=8980 $Y=52750 $D=111
M7864 157 3271 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-13 $X=9470 $Y=51990 $D=111
M7865 VDD 797 3272 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=10580 $Y=52750 $D=111
M7866 183 3272 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=11070 $Y=51990 $D=111
M7867 VDD 318 3273 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=86580 $Y=23950 $D=111
M7868 300 3273 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=87070 $Y=23190 $D=111
M7869 VDD 306 3274 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=88180 $Y=23950 $D=111
M7870 345 3274 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=88670 $Y=23190 $D=111
M7871 VDD 377 3275 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=92980 $Y=21110 $D=111
M7872 318 3275 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=93470 $Y=21110 $D=111
M7873 VDD 345 3276 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=94580 $Y=21110 $D=111
M7874 368 3276 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=95070 $Y=21110 $D=111
M7875 VDD 329 3277 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=98580 $Y=28310 $D=111
M7876 407 3277 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=99070 $Y=28310 $D=111
M7877 VDD 377 3278 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=100180 $Y=28310 $D=111
M7878 409 3278 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=100670 $Y=28310 $D=111
M7879 VDD 377 3279 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=102980 $Y=21110 $D=111
M7880 399 3279 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=103470 $Y=21110 $D=111
M7881 VDD 368 3280 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=104580 $Y=21110 $D=111
M7882 396 3280 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=105070 $Y=21110 $D=111
M7883 VDD 390 3281 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=106180 $Y=21110 $D=111
M7884 data_out[0] 3281 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=106670 $Y=21110 $D=111
M7885 VDD 399 3282 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=107780 $Y=21110 $D=111
M7886 408 3282 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=108270 $Y=21110 $D=111
M7887 VDD 543 3283 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=141780 $Y=49910 $D=111
M7888 544 3283 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=142270 $Y=49910 $D=111
M7889 VDD 544 3284 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=143380 $Y=49910 $D=111
M7890 697 3284 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=143870 $Y=49910 $D=111
M7891 VDD 611 3285 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=153380 $Y=21110 $D=111
M7892 682 3285 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=153870 $Y=21110 $D=111
M7893 VDD 570 3286 VDD lppfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16628e-13 as=2.16e-13 pd=9.80217e-07 ps=1.88e-06 nrd=0.39996 nrs=0.740741 sa=4e-07 sb=8.1e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=4.8e-15 panw9=0 panw10=0 $X=154980 $Y=21110 $D=111
M7894 620 3286 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.16e-13 as=2.80772e-13 pd=3.24e-06 ps=2.35978e-06 nrd=0.246154 nrs=0.166137 sa=5.21692e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=155470 $Y=21110 $D=111
M7895 3297 97 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=11660 $Y=9080 $D=111
M7896 3290 3292 3297 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=11980 $Y=9080 $D=111
M7897 VDD 76 3290 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=12460 $Y=9080 $D=111
M7898 VDD clk 3289 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=12980 $Y=9670 $D=111
M7899 3292 3289 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=13490 $Y=9770 $D=111
M7900 3299 3289 3290 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=14050 $Y=9310 $D=111
M7901 VDD 3291 3299 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=14370 $Y=9310 $D=111
M7902 3291 3290 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=14910 $Y=9310 $D=111
M7903 3293 3289 3291 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=15740 $Y=9060 $D=111
M7904 3302 3292 3293 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=16470 $Y=9060 $D=111
M7905 VDD 3295 3302 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=16800 $Y=9060 $D=111
M7906 3295 76 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=17260 $Y=9130 $D=111
M7907 VDD 3293 3295 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=17820 $Y=8840 $D=111
M7908 3294 3295 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=18430 $Y=9480 $D=111
M7909 VDD 3294 3287 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=19370 $Y=9610 $D=111
M7910 weight_out[0] 3295 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=19870 $Y=9610 $D=111
M7911 3313 79 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=20860 $Y=9080 $D=111
M7912 3306 3308 3313 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=21180 $Y=9080 $D=111
M7913 VDD 76 3306 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=21660 $Y=9080 $D=111
M7914 VDD clk 3305 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=22180 $Y=9670 $D=111
M7915 3308 3305 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=22690 $Y=9770 $D=111
M7916 3315 3305 3306 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=23250 $Y=9310 $D=111
M7917 VDD 3307 3315 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=23570 $Y=9310 $D=111
M7918 3307 3306 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=24110 $Y=9310 $D=111
M7919 3309 3305 3307 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=24940 $Y=9060 $D=111
M7920 3318 3308 3309 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=25670 $Y=9060 $D=111
M7921 VDD 3311 3318 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=26000 $Y=9060 $D=111
M7922 3311 76 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=26460 $Y=9130 $D=111
M7923 VDD 3309 3311 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=27020 $Y=8840 $D=111
M7924 3310 3311 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=27630 $Y=9480 $D=111
M7925 VDD 3310 3288 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=28570 $Y=9610 $D=111
M7926 weight_out[2] 3311 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=29070 $Y=9610 $D=111
M7927 3331 113 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=30060 $Y=9080 $D=111
M7928 3324 3326 3331 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=30380 $Y=9080 $D=111
M7929 VDD 128 3324 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=30860 $Y=9080 $D=111
M7930 VDD clk 3323 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=31380 $Y=9670 $D=111
M7931 3326 3323 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=31890 $Y=9770 $D=111
M7932 3333 3323 3324 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=32450 $Y=9310 $D=111
M7933 VDD 3325 3333 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=32770 $Y=9310 $D=111
M7934 3325 3324 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=33310 $Y=9310 $D=111
M7935 3327 3323 3325 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=34140 $Y=9060 $D=111
M7936 3336 3326 3327 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=34870 $Y=9060 $D=111
M7937 VDD 3329 3336 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=35200 $Y=9060 $D=111
M7938 3329 128 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=35660 $Y=9130 $D=111
M7939 VDD 3327 3329 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=36220 $Y=8840 $D=111
M7940 3328 3329 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=36830 $Y=9480 $D=111
M7941 VDD 3328 3321 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=37770 $Y=9610 $D=111
M7942 weight_out[1] 3329 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=38270 $Y=9610 $D=111
M7943 3347 195 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=39260 $Y=9080 $D=111
M7944 3340 3342 3347 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=39580 $Y=9080 $D=111
M7945 VDD 202 3340 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=40060 $Y=9080 $D=111
M7946 VDD clk 3339 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=40580 $Y=9670 $D=111
M7947 3342 3339 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=41090 $Y=9770 $D=111
M7948 3349 3339 3340 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=41650 $Y=9310 $D=111
M7949 VDD 3341 3349 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=41970 $Y=9310 $D=111
M7950 3341 3340 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=42510 $Y=9310 $D=111
M7951 3343 3339 3341 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=43340 $Y=9060 $D=111
M7952 3352 3342 3343 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=44070 $Y=9060 $D=111
M7953 VDD 3345 3352 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=44400 $Y=9060 $D=111
M7954 3345 202 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=44860 $Y=9130 $D=111
M7955 VDD 3343 3345 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=45420 $Y=8840 $D=111
M7956 3344 3345 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=46030 $Y=9480 $D=111
M7957 VDD 3344 3322 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=46970 $Y=9610 $D=111
M7958 weight_out[6] 3345 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=47470 $Y=9610 $D=111
M7959 3365 135 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=36060 $Y=14640 $D=111
M7960 3358 3360 3365 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=36380 $Y=14640 $D=111
M7961 VDD 128 3358 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=36860 $Y=14640 $D=111
M7962 VDD clk 3357 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=37380 $Y=13910 $D=111
M7963 3360 3357 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=37890 $Y=13950 $D=111
M7964 3367 3357 3358 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=38450 $Y=14410 $D=111
M7965 VDD 3359 3367 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=38770 $Y=14410 $D=111
M7966 3359 3358 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=39310 $Y=14410 $D=111
M7967 3361 3357 3359 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=40140 $Y=14660 $D=111
M7968 3370 3360 3361 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=40870 $Y=14660 $D=111
M7969 VDD 3363 3370 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=41200 $Y=14660 $D=111
M7970 3363 128 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=41660 $Y=14590 $D=111
M7971 VDD 3361 3363 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=42220 $Y=14880 $D=111
M7972 3362 3363 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=42830 $Y=14240 $D=111
M7973 VDD 3362 3355 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=43770 $Y=14050 $D=111
M7974 weight_out[4] 3363 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=44270 $Y=14050 $D=111
M7975 3381 170 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=45260 $Y=14640 $D=111
M7976 3374 3376 3381 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=45580 $Y=14640 $D=111
M7977 VDD 128 3374 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=46060 $Y=14640 $D=111
M7978 VDD clk 3373 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=46580 $Y=13910 $D=111
M7979 3376 3373 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=47090 $Y=13950 $D=111
M7980 3383 3373 3374 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=47650 $Y=14410 $D=111
M7981 VDD 3375 3383 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=47970 $Y=14410 $D=111
M7982 3375 3374 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=48510 $Y=14410 $D=111
M7983 3377 3373 3375 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=49340 $Y=14660 $D=111
M7984 3386 3376 3377 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=50070 $Y=14660 $D=111
M7985 VDD 3379 3386 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=50400 $Y=14660 $D=111
M7986 3379 128 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=50860 $Y=14590 $D=111
M7987 VDD 3377 3379 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=51420 $Y=14880 $D=111
M7988 3378 3379 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=52030 $Y=14240 $D=111
M7989 VDD 3378 3356 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=52970 $Y=14050 $D=111
M7990 weight_out[5] 3379 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=53470 $Y=14050 $D=111
M7991 3399 240 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=50460 $Y=9080 $D=111
M7992 3392 3394 3399 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=50780 $Y=9080 $D=111
M7993 VDD 202 3392 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=51260 $Y=9080 $D=111
M7994 VDD clk 3391 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=51780 $Y=9670 $D=111
M7995 3394 3391 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=52290 $Y=9770 $D=111
M7996 3401 3391 3392 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=52850 $Y=9310 $D=111
M7997 VDD 3393 3401 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=53170 $Y=9310 $D=111
M7998 3393 3392 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=53710 $Y=9310 $D=111
M7999 3395 3391 3393 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=54540 $Y=9060 $D=111
M8000 3404 3394 3395 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=55270 $Y=9060 $D=111
M8001 VDD 3397 3404 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=55600 $Y=9060 $D=111
M8002 3397 202 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=56060 $Y=9130 $D=111
M8003 VDD 3395 3397 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=56620 $Y=8840 $D=111
M8004 3396 3397 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=57230 $Y=9480 $D=111
M8005 VDD 3396 3389 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=58170 $Y=9610 $D=111
M8006 weight_out[7] 3397 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=58670 $Y=9610 $D=111
M8007 3415 310 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=59660 $Y=9080 $D=111
M8008 3408 3410 3415 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=59980 $Y=9080 $D=111
M8009 VDD 252 3408 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=60460 $Y=9080 $D=111
M8010 VDD clk 3407 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=60980 $Y=9670 $D=111
M8011 3410 3407 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=61490 $Y=9770 $D=111
M8012 3417 3407 3408 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=62050 $Y=9310 $D=111
M8013 VDD 3409 3417 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=62370 $Y=9310 $D=111
M8014 3409 3408 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=62910 $Y=9310 $D=111
M8015 3411 3407 3409 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=63740 $Y=9060 $D=111
M8016 3420 3410 3411 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=64470 $Y=9060 $D=111
M8017 VDD 3413 3420 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=64800 $Y=9060 $D=111
M8018 3413 252 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=65260 $Y=9130 $D=111
M8019 VDD 3411 3413 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=65820 $Y=8840 $D=111
M8020 3412 3413 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=66430 $Y=9480 $D=111
M8021 VDD 3412 3390 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=67370 $Y=9610 $D=111
M8022 fire_out 3413 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=67870 $Y=9610 $D=111
M8023 3433 251 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=68860 $Y=9080 $D=111
M8024 3426 3428 3433 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=69180 $Y=9080 $D=111
M8025 VDD 252 3426 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=69660 $Y=9080 $D=111
M8026 VDD clk 3425 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=70180 $Y=9670 $D=111
M8027 3428 3425 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=70690 $Y=9770 $D=111
M8028 3435 3425 3426 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=71250 $Y=9310 $D=111
M8029 VDD 3427 3435 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=71570 $Y=9310 $D=111
M8030 3427 3426 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=72110 $Y=9310 $D=111
M8031 3429 3425 3427 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=72940 $Y=9060 $D=111
M8032 3438 3428 3429 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=73670 $Y=9060 $D=111
M8033 VDD 3431 3438 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=74000 $Y=9060 $D=111
M8034 3431 252 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=74460 $Y=9130 $D=111
M8035 VDD 3429 3431 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=75020 $Y=8840 $D=111
M8036 3430 3431 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=75630 $Y=9480 $D=111
M8037 VDD 3430 3423 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=76570 $Y=9610 $D=111
M8038 result[1] 3431 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=77070 $Y=9610 $D=111
M8039 3449 828 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=78060 $Y=9080 $D=111
M8040 3442 3444 3449 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=78380 $Y=9080 $D=111
M8041 VDD 299 3442 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=78860 $Y=9080 $D=111
M8042 VDD clk 3441 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=79380 $Y=9670 $D=111
M8043 3444 3441 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=79890 $Y=9770 $D=111
M8044 3451 3441 3442 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=80450 $Y=9310 $D=111
M8045 VDD 3443 3451 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=80770 $Y=9310 $D=111
M8046 3443 3442 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=81310 $Y=9310 $D=111
M8047 3445 3441 3443 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=82140 $Y=9060 $D=111
M8048 3454 3444 3445 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=82870 $Y=9060 $D=111
M8049 VDD 3447 3454 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=83200 $Y=9060 $D=111
M8050 3447 299 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=83660 $Y=9130 $D=111
M8051 VDD 3445 3447 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=84220 $Y=8840 $D=111
M8052 3446 3447 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=84830 $Y=9480 $D=111
M8053 VDD 3446 3424 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=85770 $Y=9610 $D=111
M8054 result[2] 3447 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=86270 $Y=9610 $D=111
M8055 3467 305 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=80060 $Y=29040 $D=111
M8056 3460 3462 3467 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=80380 $Y=29040 $D=111
M8057 VDD 303 3460 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=80860 $Y=29040 $D=111
M8058 VDD clk 3459 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=81380 $Y=28310 $D=111
M8059 3462 3459 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=81890 $Y=28350 $D=111
M8060 3469 3459 3460 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=82450 $Y=28810 $D=111
M8061 VDD 3461 3469 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=82770 $Y=28810 $D=111
M8062 3461 3460 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=83310 $Y=28810 $D=111
M8063 3463 3459 3461 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=84140 $Y=29060 $D=111
M8064 3472 3462 3463 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=84870 $Y=29060 $D=111
M8065 VDD 3465 3472 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=85200 $Y=29060 $D=111
M8066 3465 303 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=85660 $Y=28990 $D=111
M8067 VDD 3463 3465 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=86220 $Y=29280 $D=111
M8068 3464 3465 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=86830 $Y=28640 $D=111
M8069 VDD 3464 3457 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=87770 $Y=28450 $D=111
M8070 result[5] 3465 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=88270 $Y=28450 $D=111
M8071 3483 217 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=89260 $Y=29040 $D=111
M8072 3476 3478 3483 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=89580 $Y=29040 $D=111
M8073 VDD 329 3476 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=90060 $Y=29040 $D=111
M8074 VDD clk 3475 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=90580 $Y=28310 $D=111
M8075 3478 3475 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=91090 $Y=28350 $D=111
M8076 3485 3475 3476 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=91650 $Y=28810 $D=111
M8077 VDD 3477 3485 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=91970 $Y=28810 $D=111
M8078 3477 3476 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=92510 $Y=28810 $D=111
M8079 3479 3475 3477 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=93340 $Y=29060 $D=111
M8080 3488 3478 3479 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=94070 $Y=29060 $D=111
M8081 VDD 3481 3488 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=94400 $Y=29060 $D=111
M8082 3481 329 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=94860 $Y=28990 $D=111
M8083 VDD 3479 3481 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=95420 $Y=29280 $D=111
M8084 3480 3481 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=96030 $Y=28640 $D=111
M8085 VDD 3480 3458 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=96970 $Y=28450 $D=111
M8086 390 3481 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=97470 $Y=28450 $D=111
M8087 3501 333 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=87260 $Y=9080 $D=111
M8088 3494 3496 3501 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=87580 $Y=9080 $D=111
M8089 VDD 356 3494 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=88060 $Y=9080 $D=111
M8090 VDD clk 3493 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=88580 $Y=9670 $D=111
M8091 3496 3493 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=89090 $Y=9770 $D=111
M8092 3503 3493 3494 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=89650 $Y=9310 $D=111
M8093 VDD 3495 3503 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=89970 $Y=9310 $D=111
M8094 3495 3494 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=90510 $Y=9310 $D=111
M8095 3497 3493 3495 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=91340 $Y=9060 $D=111
M8096 3506 3496 3497 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=92070 $Y=9060 $D=111
M8097 VDD 3499 3506 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=92400 $Y=9060 $D=111
M8098 3499 356 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=92860 $Y=9130 $D=111
M8099 VDD 3497 3499 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=93420 $Y=8840 $D=111
M8100 3498 3499 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=94030 $Y=9480 $D=111
M8101 VDD 3498 3491 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=94970 $Y=9610 $D=111
M8102 result[3] 3499 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=95470 $Y=9610 $D=111
M8103 3517 364 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=96460 $Y=9080 $D=111
M8104 3510 3512 3517 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=96780 $Y=9080 $D=111
M8105 VDD 356 3510 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=97260 $Y=9080 $D=111
M8106 VDD clk 3509 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=97780 $Y=9670 $D=111
M8107 3512 3509 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=98290 $Y=9770 $D=111
M8108 3519 3509 3510 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=98850 $Y=9310 $D=111
M8109 VDD 3511 3519 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=99170 $Y=9310 $D=111
M8110 3511 3510 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=99710 $Y=9310 $D=111
M8111 3513 3509 3511 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=100540 $Y=9060 $D=111
M8112 3522 3512 3513 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=101270 $Y=9060 $D=111
M8113 VDD 3515 3522 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=101600 $Y=9060 $D=111
M8114 3515 356 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=102060 $Y=9130 $D=111
M8115 VDD 3513 3515 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=102620 $Y=8840 $D=111
M8116 3514 3515 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=103230 $Y=9480 $D=111
M8117 VDD 3514 3492 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=104170 $Y=9610 $D=111
M8118 result[10] 3515 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=104670 $Y=9610 $D=111
M8119 3535 332 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=89660 $Y=23480 $D=111
M8120 3528 3530 3535 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=89980 $Y=23480 $D=111
M8121 VDD 329 3528 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=90460 $Y=23480 $D=111
M8122 VDD clk 3527 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=90980 $Y=24070 $D=111
M8123 3530 3527 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=91490 $Y=24170 $D=111
M8124 3537 3527 3528 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=92050 $Y=23710 $D=111
M8125 VDD 3529 3537 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=92370 $Y=23710 $D=111
M8126 3529 3528 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=92910 $Y=23710 $D=111
M8127 3531 3527 3529 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=93740 $Y=23460 $D=111
M8128 3540 3530 3531 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=94470 $Y=23460 $D=111
M8129 VDD 3533 3540 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=94800 $Y=23460 $D=111
M8130 3533 329 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=95260 $Y=23530 $D=111
M8131 VDD 3531 3533 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=95820 $Y=23240 $D=111
M8132 3532 3533 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=96430 $Y=23880 $D=111
M8133 VDD 3532 3525 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=97370 $Y=24010 $D=111
M8134 result[7] 3533 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=97870 $Y=24010 $D=111
M8135 3551 832 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=98860 $Y=23480 $D=111
M8136 3544 3546 3551 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=99180 $Y=23480 $D=111
M8137 VDD 407 3544 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=99660 $Y=23480 $D=111
M8138 VDD clk 3543 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=100180 $Y=24070 $D=111
M8139 3546 3543 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=100690 $Y=24170 $D=111
M8140 3553 3543 3544 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=101250 $Y=23710 $D=111
M8141 VDD 3545 3553 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=101570 $Y=23710 $D=111
M8142 3545 3544 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=102110 $Y=23710 $D=111
M8143 3547 3543 3545 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=102940 $Y=23460 $D=111
M8144 3556 3546 3547 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=103670 $Y=23460 $D=111
M8145 VDD 3549 3556 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=104000 $Y=23460 $D=111
M8146 3549 407 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=104460 $Y=23530 $D=111
M8147 VDD 3547 3549 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=105020 $Y=23240 $D=111
M8148 3548 3549 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=105630 $Y=23880 $D=111
M8149 VDD 3548 3526 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=106570 $Y=24010 $D=111
M8150 result[8] 3549 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=107070 $Y=24010 $D=111
M8151 3569 388 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=105260 $Y=14640 $D=111
M8152 3562 3564 3569 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=105580 $Y=14640 $D=111
M8153 VDD 371 3562 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=106060 $Y=14640 $D=111
M8154 VDD clk 3561 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=106580 $Y=13910 $D=111
M8155 3564 3561 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=107090 $Y=13950 $D=111
M8156 3571 3561 3562 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=107650 $Y=14410 $D=111
M8157 VDD 3563 3571 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=107970 $Y=14410 $D=111
M8158 3563 3562 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=108510 $Y=14410 $D=111
M8159 3565 3561 3563 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=109340 $Y=14660 $D=111
M8160 3574 3564 3565 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=110070 $Y=14660 $D=111
M8161 VDD 3567 3574 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=110400 $Y=14660 $D=111
M8162 3567 371 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=110860 $Y=14590 $D=111
M8163 VDD 3565 3567 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=111420 $Y=14880 $D=111
M8164 3566 3567 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=112030 $Y=14240 $D=111
M8165 VDD 3566 3559 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=112970 $Y=14050 $D=111
M8166 result[12] 3567 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=113470 $Y=14050 $D=111
M8167 3585 424 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=114460 $Y=14640 $D=111
M8168 3578 3580 3585 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=114780 $Y=14640 $D=111
M8169 VDD 428 3578 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=115260 $Y=14640 $D=111
M8170 VDD clk 3577 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=115780 $Y=13910 $D=111
M8171 3580 3577 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=116290 $Y=13950 $D=111
M8172 3587 3577 3578 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=116850 $Y=14410 $D=111
M8173 VDD 3579 3587 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=117170 $Y=14410 $D=111
M8174 3579 3578 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=117710 $Y=14410 $D=111
M8175 3581 3577 3579 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=118540 $Y=14660 $D=111
M8176 3590 3580 3581 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=119270 $Y=14660 $D=111
M8177 VDD 3583 3590 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=119600 $Y=14660 $D=111
M8178 3583 428 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=120060 $Y=14590 $D=111
M8179 VDD 3581 3583 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=120620 $Y=14880 $D=111
M8180 3582 3583 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=121230 $Y=14240 $D=111
M8181 VDD 3582 3560 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=122170 $Y=14050 $D=111
M8182 result[15] 3583 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=122670 $Y=14050 $D=111
M8183 3603 449 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=119260 $Y=9080 $D=111
M8184 3596 3598 3603 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=119580 $Y=9080 $D=111
M8185 VDD 479 3596 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=120060 $Y=9080 $D=111
M8186 VDD clk 3595 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=120580 $Y=9670 $D=111
M8187 3598 3595 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=121090 $Y=9770 $D=111
M8188 3605 3595 3596 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=121650 $Y=9310 $D=111
M8189 VDD 3597 3605 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=121970 $Y=9310 $D=111
M8190 3597 3596 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=122510 $Y=9310 $D=111
M8191 3599 3595 3597 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=123340 $Y=9060 $D=111
M8192 3608 3598 3599 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=124070 $Y=9060 $D=111
M8193 VDD 3601 3608 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=124400 $Y=9060 $D=111
M8194 3601 479 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=124860 $Y=9130 $D=111
M8195 VDD 3599 3601 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=125420 $Y=8840 $D=111
M8196 3600 3601 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=126030 $Y=9480 $D=111
M8197 VDD 3600 3593 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=126970 $Y=9610 $D=111
M8198 result[16] 3601 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=127470 $Y=9610 $D=111
M8199 3619 513 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=128460 $Y=9080 $D=111
M8200 3612 3614 3619 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=128780 $Y=9080 $D=111
M8201 VDD 479 3612 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=129260 $Y=9080 $D=111
M8202 VDD clk 3611 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=129780 $Y=9670 $D=111
M8203 3614 3611 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=130290 $Y=9770 $D=111
M8204 3621 3611 3612 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=130850 $Y=9310 $D=111
M8205 VDD 3613 3621 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=131170 $Y=9310 $D=111
M8206 3613 3612 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=131710 $Y=9310 $D=111
M8207 3615 3611 3613 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=132540 $Y=9060 $D=111
M8208 3624 3614 3615 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=133270 $Y=9060 $D=111
M8209 VDD 3617 3624 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=133600 $Y=9060 $D=111
M8210 3617 479 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=134060 $Y=9130 $D=111
M8211 VDD 3615 3617 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=134620 $Y=8840 $D=111
M8212 3616 3617 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=135230 $Y=9480 $D=111
M8213 VDD 3616 3594 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=136170 $Y=9610 $D=111
M8214 result[17] 3617 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=136670 $Y=9610 $D=111
M8215 3637 541 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=137660 $Y=9080 $D=111
M8216 3630 3632 3637 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=137980 $Y=9080 $D=111
M8217 VDD 584 3630 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=138460 $Y=9080 $D=111
M8218 VDD clk 3629 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=138980 $Y=9670 $D=111
M8219 3632 3629 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=139490 $Y=9770 $D=111
M8220 3639 3629 3630 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=140050 $Y=9310 $D=111
M8221 VDD 3631 3639 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=140370 $Y=9310 $D=111
M8222 3631 3630 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=140910 $Y=9310 $D=111
M8223 3633 3629 3631 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=141740 $Y=9060 $D=111
M8224 3642 3632 3633 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=142470 $Y=9060 $D=111
M8225 VDD 3635 3642 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=142800 $Y=9060 $D=111
M8226 3635 584 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=143260 $Y=9130 $D=111
M8227 VDD 3633 3635 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=143820 $Y=8840 $D=111
M8228 3634 3635 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=144430 $Y=9480 $D=111
M8229 VDD 3634 3627 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=145370 $Y=9610 $D=111
M8230 result[18] 3635 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=145870 $Y=9610 $D=111
M8231 3653 604 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=146860 $Y=9080 $D=111
M8232 3646 3648 3653 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=147180 $Y=9080 $D=111
M8233 VDD 584 3646 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=147660 $Y=9080 $D=111
M8234 VDD clk 3645 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=3.96e-14 $X=148180 $Y=9670 $D=111
M8235 3648 3645 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=2.76e-14 $X=148690 $Y=9770 $D=111
M8236 3655 3645 3646 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=149250 $Y=9310 $D=111
M8237 VDD 3647 3655 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=149570 $Y=9310 $D=111
M8238 3647 3646 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=2.04e-14 panw10=2.28e-14 $X=150110 $Y=9310 $D=111
M8239 3649 3645 3647 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=150940 $Y=9060 $D=111
M8240 3658 3648 3649 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=151670 $Y=9060 $D=111
M8241 VDD 3651 3658 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=6.72e-14 panw10=0 $X=152000 $Y=9060 $D=111
M8242 3651 584 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=6.36e-14 panw10=1.2e-15 $X=152460 $Y=9130 $D=111
M8243 VDD 3649 3651 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=3e-14 panw10=1.8e-14 $X=153020 $Y=8840 $D=111
M8244 3650 3651 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=3.36e-14 $X=153630 $Y=9480 $D=111
M8245 VDD 3650 3628 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=154570 $Y=9610 $D=111
M8246 result[21] 3651 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=4.08e-14 $X=155070 $Y=9610 $D=111
M8247 3671 579 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=140860 $Y=14640 $D=111
M8248 3664 3666 3671 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=141180 $Y=14640 $D=111
M8249 VDD 584 3664 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=141660 $Y=14640 $D=111
M8250 VDD clk 3663 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=142180 $Y=13910 $D=111
M8251 3666 3663 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=142690 $Y=13950 $D=111
M8252 3673 3663 3664 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=143250 $Y=14410 $D=111
M8253 VDD 3665 3673 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=143570 $Y=14410 $D=111
M8254 3665 3664 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=144110 $Y=14410 $D=111
M8255 3667 3663 3665 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=144940 $Y=14660 $D=111
M8256 3676 3666 3667 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=145670 $Y=14660 $D=111
M8257 VDD 3669 3676 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=146000 $Y=14660 $D=111
M8258 3669 584 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=146460 $Y=14590 $D=111
M8259 VDD 3667 3669 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=147020 $Y=14880 $D=111
M8260 3668 3669 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=147630 $Y=14240 $D=111
M8261 VDD 3668 3661 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=148570 $Y=14050 $D=111
M8262 result[19] 3669 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=149070 $Y=14050 $D=111
M8263 3687 623 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=150060 $Y=14640 $D=111
M8264 3680 3682 3687 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=150380 $Y=14640 $D=111
M8265 VDD 638 3680 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=150860 $Y=14640 $D=111
M8266 VDD clk 3679 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=151380 $Y=13910 $D=111
M8267 3682 3679 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=151890 $Y=13950 $D=111
M8268 3689 3679 3680 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=152450 $Y=14410 $D=111
M8269 VDD 3681 3689 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=152770 $Y=14410 $D=111
M8270 3681 3680 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=153310 $Y=14410 $D=111
M8271 3683 3679 3681 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=154140 $Y=14660 $D=111
M8272 3692 3682 3683 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=154870 $Y=14660 $D=111
M8273 VDD 3685 3692 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=155200 $Y=14660 $D=111
M8274 3685 638 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=155660 $Y=14590 $D=111
M8275 VDD 3683 3685 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=156220 $Y=14880 $D=111
M8276 3684 3685 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=156830 $Y=14240 $D=111
M8277 VDD 3684 3662 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=157770 $Y=14050 $D=111
M8278 result[20] 3685 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=158270 $Y=14050 $D=111
M8279 3705 612 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=149260 $Y=29040 $D=111
M8280 3698 3700 3705 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=149580 $Y=29040 $D=111
M8281 VDD 662 3698 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=150060 $Y=29040 $D=111
M8282 VDD clk 3697 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=150580 $Y=28310 $D=111
M8283 3700 3697 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=151090 $Y=28350 $D=111
M8284 3707 3697 3698 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=151650 $Y=28810 $D=111
M8285 VDD 3699 3707 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=151970 $Y=28810 $D=111
M8286 3699 3698 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=152510 $Y=28810 $D=111
M8287 3701 3697 3699 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=153340 $Y=29060 $D=111
M8288 3710 3700 3701 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=154070 $Y=29060 $D=111
M8289 VDD 3703 3710 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=154400 $Y=29060 $D=111
M8290 3703 662 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=154860 $Y=28990 $D=111
M8291 VDD 3701 3703 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=155420 $Y=29280 $D=111
M8292 3702 3703 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=156030 $Y=28640 $D=111
M8293 VDD 3702 3695 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=156970 $Y=28450 $D=111
M8294 result[25] 3703 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=157470 $Y=28450 $D=111
M8295 3721 656 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=158460 $Y=29040 $D=111
M8296 3714 3716 3721 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=158780 $Y=29040 $D=111
M8297 VDD 641 3714 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=159260 $Y=29040 $D=111
M8298 VDD clk 3713 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=159780 $Y=28310 $D=111
M8299 3716 3713 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-15 panw8=0 panw9=0 panw10=0 $X=160290 $Y=28350 $D=111
M8300 3723 3713 3714 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=160850 $Y=28810 $D=111
M8301 VDD 3715 3723 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=161170 $Y=28810 $D=111
M8302 3715 3714 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=161710 $Y=28810 $D=111
M8303 3717 3713 3715 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=162540 $Y=29060 $D=111
M8304 3726 3716 3717 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=163270 $Y=29060 $D=111
M8305 VDD 3719 3726 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=163600 $Y=29060 $D=111
M8306 3719 641 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=164060 $Y=28990 $D=111
M8307 VDD 3717 3719 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3343e-13 as=8.48e-14 pd=9.32598e-07 ps=1.01e-06 nrd=1.70191 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=164620 $Y=29280 $D=111
M8308 3718 3719 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.3343e-13 pd=1.2e-06 ps=9.32598e-07 nrd=1.14286 nrs=1.70191 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=165230 $Y=28640 $D=111
M8309 VDD 3718 3696 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62022e-13 as=1.088e-13 pd=1.13244e-06 ps=1.32e-06 nrd=1.40157 nrs=0.941176 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=166170 $Y=28450 $D=111
M8310 result[26] 3719 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.088e-13 as=1.62022e-13 pd=1.32e-06 ps=1.13244e-06 nrd=0.941176 nrs=1.40157 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.16e-14 panw8=0 panw9=0 panw10=0 $X=166670 $Y=28450 $D=111
M8311 VDD 228 3729 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.91478e-14 as=9.24e-14 pd=6.33043e-07 ps=1.22e-06 nrd=0.881988 nrs=1.17857 sa=3.3e-07 sb=1.37e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.32e-14 panw8=0 panw9=0 panw10=0 $X=61620 $Y=52880 $D=111
M8312 221 241 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.58052e-13 pd=1e-06 ps=1.44696e-06 nrd=0.28125 nrs=0.38587 sa=5.51875e-07 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=62140 $Y=52520 $D=111
M8313 VDD 3729 221 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.267e-13 as=1.152e-13 pd=2.64e-06 ps=1e-06 nrd=0.797607 nrs=0.28125 sa=1.03187e-06 sb=3.7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=62620 $Y=52520 $D=111
M8314 VDD 437 3731 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.91478e-14 as=9.24e-14 pd=6.33043e-07 ps=1.22e-06 nrd=0.881988 nrs=1.17857 sa=3.3e-07 sb=1.37e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.32e-14 panw8=0 panw9=0 panw10=0 $X=112420 $Y=57240 $D=111
M8315 412 430 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.58052e-13 pd=1e-06 ps=1.44696e-06 nrd=0.28125 nrs=0.38587 sa=5.51875e-07 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=112940 $Y=57240 $D=111
M8316 VDD 3731 412 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.267e-13 as=1.152e-13 pd=2.64e-06 ps=1e-06 nrd=0.797607 nrs=0.28125 sa=1.03187e-06 sb=3.7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=113420 $Y=57240 $D=111
M8317 VDD 562 3733 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.91478e-14 as=9.24e-14 pd=6.33043e-07 ps=1.22e-06 nrd=0.881988 nrs=1.17857 sa=3.3e-07 sb=1.37e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.32e-14 panw8=0 panw9=0 panw10=0 $X=138020 $Y=67280 $D=111
M8318 913 539 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.58052e-13 pd=1e-06 ps=1.44696e-06 nrd=0.28125 nrs=0.38587 sa=5.51875e-07 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=138540 $Y=66920 $D=111
M8319 VDD 3733 913 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.267e-13 as=1.152e-13 pd=2.64e-06 ps=1e-06 nrd=0.797607 nrs=0.28125 sa=1.03187e-06 sb=3.7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=139020 $Y=66920 $D=111
M8320 VDD 559 3735 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.91478e-14 as=9.24e-14 pd=6.33043e-07 ps=1.22e-06 nrd=0.881988 nrs=1.17857 sa=3.3e-07 sb=1.37e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.32e-14 panw8=0 panw9=0 panw10=0 $X=138420 $Y=60080 $D=111
M8321 553 549 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.58052e-13 pd=1e-06 ps=1.44696e-06 nrd=0.28125 nrs=0.38587 sa=5.51875e-07 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=138940 $Y=59720 $D=111
M8322 VDD 3735 553 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.267e-13 as=1.152e-13 pd=2.64e-06 ps=1e-06 nrd=0.797607 nrs=0.28125 sa=1.03187e-06 sb=3.7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=139420 $Y=59720 $D=111
M8323 VDD 575 3737 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.91478e-14 as=9.24e-14 pd=6.33043e-07 ps=1.22e-06 nrd=0.881988 nrs=1.17857 sa=3.3e-07 sb=1.37e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.32e-14 panw8=0 panw9=0 panw10=0 $X=143620 $Y=60080 $D=111
M8324 567 560 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.58052e-13 pd=1e-06 ps=1.44696e-06 nrd=0.28125 nrs=0.38587 sa=5.51875e-07 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=144140 $Y=59720 $D=111
M8325 VDD 3737 567 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.267e-13 as=1.152e-13 pd=2.64e-06 ps=1e-06 nrd=0.797607 nrs=0.28125 sa=1.03187e-06 sb=3.7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=2.4e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=144620 $Y=59720 $D=111
M8326 87 82 VDD VDD lppfet w=1.24e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.29877e-13 as=3.968e-13 pd=1.69573e-06 ps=3.12e-06 nrd=0.149504 nrs=0.258065 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=26810 $Y=57160 $D=111
M8327 VDD 82 87 VDD lppfet w=1.1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.48643e-13 as=2.03923e-13 pd=3.00143e-06 ps=1.50427e-06 nrd=0.370779 nrs=0.168531 sa=8e-07 sb=4.1e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=27290 $Y=57160 $D=111
M8328 148 97 VDD VDD lppfet w=1.24e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.29877e-13 as=3.968e-13 pd=1.69573e-06 ps=3.12e-06 nrd=0.149504 nrs=0.258065 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=40810 $Y=23200 $D=111
M8329 VDD 97 148 VDD lppfet w=1.1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.48643e-13 as=2.03923e-13 pd=3.00143e-06 ps=1.50427e-06 nrd=0.370779 nrs=0.168531 sa=8e-07 sb=4.1e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=41290 $Y=23340 $D=111
M8330 411 402 VDD VDD lppfet w=1.24e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.29877e-13 as=3.968e-13 pd=1.69573e-06 ps=3.12e-06 nrd=0.149504 nrs=0.258065 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=108010 $Y=73600 $D=111
M8331 VDD 402 411 VDD lppfet w=1.1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.48643e-13 as=2.03923e-13 pd=3.00143e-06 ps=1.50427e-06 nrd=0.370779 nrs=0.168531 sa=8e-07 sb=4.1e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=108490 $Y=73740 $D=111
M8332 435 404 VDD VDD lppfet w=1.24e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.29877e-13 as=3.968e-13 pd=1.69573e-06 ps=3.12e-06 nrd=0.149504 nrs=0.258065 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=110810 $Y=71560 $D=111
M8333 VDD 404 435 VDD lppfet w=1.1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.48643e-13 as=2.03923e-13 pd=3.00143e-06 ps=1.50427e-06 nrd=0.370779 nrs=0.168531 sa=8e-07 sb=4.1e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=111290 $Y=71560 $D=111
M8334 499 523 VDD VDD lppfet w=1.24e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.29877e-13 as=3.968e-13 pd=1.69573e-06 ps=3.12e-06 nrd=0.149504 nrs=0.258065 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=133210 $Y=37600 $D=111
M8335 VDD 523 499 VDD lppfet w=1.1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.48643e-13 as=2.03923e-13 pd=3.00143e-06 ps=1.50427e-06 nrd=0.370779 nrs=0.168531 sa=8e-07 sb=4.1e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=133690 $Y=37740 $D=111
M8336 849 503 VDD VDD lppfet w=1.24e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.29877e-13 as=3.968e-13 pd=1.69573e-06 ps=3.12e-06 nrd=0.149504 nrs=0.258065 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=133610 $Y=66400 $D=111
M8337 VDD 503 849 VDD lppfet w=1.1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.48643e-13 as=2.03923e-13 pd=3.00143e-06 ps=1.50427e-06 nrd=0.370779 nrs=0.168531 sa=8e-07 sb=4.1e-07 sd=0 panw1=0 panw2=0 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=134090 $Y=66540 $D=111
M8338 3740 59 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=20810 $Y=52110 $D=111
M8339 803 63 3740 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=1.96571e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=21130 $Y=52110 $D=111
M8340 3741 63 803 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=1.82723e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=21610 $Y=52110 $D=111
M8341 VDD 59 3741 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=1.73295e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=21930 $Y=52110 $D=111
M8342 3742 59 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=1.59152e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=22410 $Y=52110 $D=111
M8343 803 63 3742 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.21737e-13 as=1.12e-13 pd=1.74222e-06 ps=1.32e-06 nrd=0.176768 nrs=0.0892857 sa=2e-06 sb=1.39848e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=22730 $Y=52110 $D=111
M8344 VDD 75 803 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55152e-13 as=1.70263e-13 pd=1.22713e-06 ps=1.33778e-06 nrd=0.209778 nrs=0.230209 sa=1.87721e-06 sb=1.36686e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=23210 $Y=52430 $D=111
M8345 803 75 VDD VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.53e-13 as=1.53348e-13 pd=1.21e-06 ps=1.21287e-06 nrd=0.211765 nrs=0.212246 sa=1.90965e-06 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=23690 $Y=52440 $D=111
M8346 VDD 75 803 VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.182e-13 as=1.53e-13 pd=2.9e-06 ps=1.21e-06 nrd=0.578824 nrs=0.211765 sa=1.94353e-06 sb=4.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=24170 $Y=52440 $D=111
M8347 3744 142 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=30010 $Y=42770 $D=111
M8348 103 84 3744 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=1.96571e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=30330 $Y=42770 $D=111
M8349 3745 84 103 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=1.82723e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=30810 $Y=42770 $D=111
M8350 VDD 142 3745 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=1.73295e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=31130 $Y=42770 $D=111
M8351 3746 142 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=1.59152e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=31610 $Y=42770 $D=111
M8352 103 84 3746 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.21737e-13 as=1.12e-13 pd=1.74222e-06 ps=1.32e-06 nrd=0.176768 nrs=0.0892857 sa=2e-06 sb=1.39848e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=31930 $Y=42770 $D=111
M8353 VDD 108 103 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55152e-13 as=1.70263e-13 pd=1.22713e-06 ps=1.33778e-06 nrd=0.209778 nrs=0.230209 sa=1.87721e-06 sb=1.36686e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=32410 $Y=42710 $D=111
M8354 103 108 VDD VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.53e-13 as=1.53348e-13 pd=1.21e-06 ps=1.21287e-06 nrd=0.211765 nrs=0.212246 sa=1.90965e-06 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=32890 $Y=42710 $D=111
M8355 VDD 108 103 VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.182e-13 as=1.53e-13 pd=2.9e-06 ps=1.21e-06 nrd=0.578824 nrs=0.211765 sa=1.94353e-06 sb=4.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=33370 $Y=42710 $D=111
M8356 3748 119 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=30410 $Y=21170 $D=111
M8357 15 118 3748 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=1.96571e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=30730 $Y=21170 $D=111
M8358 3749 118 15 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=1.82723e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=31210 $Y=21170 $D=111
M8359 VDD 119 3749 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=1.73295e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=31530 $Y=21170 $D=111
M8360 3750 119 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=1.59152e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=32010 $Y=21170 $D=111
M8361 15 118 3750 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.21737e-13 as=1.12e-13 pd=1.74222e-06 ps=1.32e-06 nrd=0.176768 nrs=0.0892857 sa=2e-06 sb=1.39848e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=32330 $Y=21170 $D=111
M8362 VDD 132 15 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55152e-13 as=1.70263e-13 pd=1.22713e-06 ps=1.33778e-06 nrd=0.209778 nrs=0.230209 sa=1.87721e-06 sb=1.36686e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=32810 $Y=21110 $D=111
M8363 15 132 VDD VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.53e-13 as=1.53348e-13 pd=1.21e-06 ps=1.21287e-06 nrd=0.211765 nrs=0.212246 sa=1.90965e-06 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=33290 $Y=21110 $D=111
M8364 VDD 132 15 VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.182e-13 as=1.53e-13 pd=2.9e-06 ps=1.21e-06 nrd=0.578824 nrs=0.211765 sa=1.94353e-06 sb=4.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=33770 $Y=21110 $D=111
M8365 3752 143 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=41610 $Y=16110 $D=111
M8366 167 177 3752 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=1.96571e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=41930 $Y=16110 $D=111
M8367 3753 177 167 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=1.82723e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=42410 $Y=16110 $D=111
M8368 VDD 143 3753 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=1.73295e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=42730 $Y=16110 $D=111
M8369 3754 143 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=1.59152e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=43210 $Y=16110 $D=111
M8370 167 177 3754 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.21737e-13 as=1.12e-13 pd=1.74222e-06 ps=1.32e-06 nrd=0.176768 nrs=0.0892857 sa=2e-06 sb=1.39848e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=43530 $Y=16110 $D=111
M8371 VDD 169 167 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55152e-13 as=1.70263e-13 pd=1.22713e-06 ps=1.33778e-06 nrd=0.209778 nrs=0.230209 sa=1.87721e-06 sb=1.36686e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=44010 $Y=16430 $D=111
M8372 167 169 VDD VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.53e-13 as=1.53348e-13 pd=1.21e-06 ps=1.21287e-06 nrd=0.211765 nrs=0.212246 sa=1.90965e-06 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=44490 $Y=16440 $D=111
M8373 VDD 169 167 VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.182e-13 as=1.53e-13 pd=2.9e-06 ps=1.21e-06 nrd=0.578824 nrs=0.211765 sa=1.94353e-06 sb=4.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=44970 $Y=16440 $D=111
M8374 3756 358 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=96010 $Y=73710 $D=111
M8375 404 353 3756 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=1.96571e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=96330 $Y=73710 $D=111
M8376 3757 353 404 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=1.82723e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=96810 $Y=73710 $D=111
M8377 VDD 358 3757 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=1.73295e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=97130 $Y=73710 $D=111
M8378 3758 358 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=1.59152e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=97610 $Y=73710 $D=111
M8379 404 353 3758 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.21737e-13 as=1.12e-13 pd=1.74222e-06 ps=1.32e-06 nrd=0.176768 nrs=0.0892857 sa=2e-06 sb=1.39848e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=97930 $Y=73710 $D=111
M8380 VDD 361 404 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55152e-13 as=1.70263e-13 pd=1.22713e-06 ps=1.33778e-06 nrd=0.209778 nrs=0.230209 sa=1.87721e-06 sb=1.36686e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=98410 $Y=74030 $D=111
M8381 404 361 VDD VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.53e-13 as=1.53348e-13 pd=1.21e-06 ps=1.21287e-06 nrd=0.211765 nrs=0.212246 sa=1.90965e-06 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=98890 $Y=74040 $D=111
M8382 VDD 361 404 VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.182e-13 as=1.53e-13 pd=2.9e-06 ps=1.21e-06 nrd=0.578824 nrs=0.211765 sa=1.94353e-06 sb=4.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=99370 $Y=74040 $D=111
M8383 3760 496 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=122410 $Y=71570 $D=111
M8384 503 402 3760 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=1.96571e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=122730 $Y=71570 $D=111
M8385 3761 402 503 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=1.82723e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=123210 $Y=71570 $D=111
M8386 VDD 496 3761 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=1.73295e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=123530 $Y=71570 $D=111
M8387 3762 496 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=1.59152e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=124010 $Y=71570 $D=111
M8388 503 402 3762 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.21737e-13 as=1.12e-13 pd=1.74222e-06 ps=1.32e-06 nrd=0.176768 nrs=0.0892857 sa=2e-06 sb=1.39848e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=124330 $Y=71570 $D=111
M8389 VDD 842 503 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55152e-13 as=1.70263e-13 pd=1.22713e-06 ps=1.33778e-06 nrd=0.209778 nrs=0.230209 sa=1.87721e-06 sb=1.36686e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=124810 $Y=71510 $D=111
M8390 503 842 VDD VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.53e-13 as=1.53348e-13 pd=1.21e-06 ps=1.21287e-06 nrd=0.211765 nrs=0.212246 sa=1.90965e-06 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=125290 $Y=71510 $D=111
M8391 VDD 842 503 VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.182e-13 as=1.53e-13 pd=2.9e-06 ps=1.21e-06 nrd=0.578824 nrs=0.211765 sa=1.94353e-06 sb=4.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=125770 $Y=71510 $D=111
M8392 3764 476 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=127210 $Y=66510 $D=111
M8393 482 846 3764 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=1.96571e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=127530 $Y=66510 $D=111
M8394 3765 846 482 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=1.82723e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=128010 $Y=66510 $D=111
M8395 VDD 476 3765 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=1.73295e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=128330 $Y=66510 $D=111
M8396 3766 476 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=1.59152e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=128810 $Y=66510 $D=111
M8397 482 846 3766 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.21737e-13 as=1.12e-13 pd=1.74222e-06 ps=1.32e-06 nrd=0.176768 nrs=0.0892857 sa=2e-06 sb=1.39848e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=129130 $Y=66510 $D=111
M8398 VDD 495 482 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55152e-13 as=1.70263e-13 pd=1.22713e-06 ps=1.33778e-06 nrd=0.209778 nrs=0.230209 sa=1.87721e-06 sb=1.36686e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=129610 $Y=66830 $D=111
M8399 482 495 VDD VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.53e-13 as=1.53348e-13 pd=1.21e-06 ps=1.21287e-06 nrd=0.211765 nrs=0.212246 sa=1.90965e-06 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=130090 $Y=66840 $D=111
M8400 VDD 495 482 VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.182e-13 as=1.53e-13 pd=2.9e-06 ps=1.21e-06 nrd=0.578824 nrs=0.211765 sa=1.94353e-06 sb=4.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=130570 $Y=66840 $D=111
M8401 3768 502 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=132810 $Y=44910 $D=111
M8402 598 512 3768 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=1.96571e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=133130 $Y=44910 $D=111
M8403 3769 512 598 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=1.82723e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=133610 $Y=44910 $D=111
M8404 VDD 502 3769 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=1.73295e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=133930 $Y=44910 $D=111
M8405 3770 502 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=1.59152e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=134410 $Y=44910 $D=111
M8406 598 512 3770 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.21737e-13 as=1.12e-13 pd=1.74222e-06 ps=1.32e-06 nrd=0.176768 nrs=0.0892857 sa=2e-06 sb=1.39848e-06 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=134730 $Y=44910 $D=111
M8407 VDD 532 598 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.55152e-13 as=1.70263e-13 pd=1.22713e-06 ps=1.33778e-06 nrd=0.209778 nrs=0.230209 sa=1.87721e-06 sb=1.36686e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=135210 $Y=45230 $D=111
M8408 598 532 VDD VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.53e-13 as=1.53348e-13 pd=1.21e-06 ps=1.21287e-06 nrd=0.211765 nrs=0.212246 sa=1.90965e-06 sb=9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=135690 $Y=45240 $D=111
M8409 VDD 532 598 VDD lppfet w=8.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.182e-13 as=1.53e-13 pd=2.9e-06 ps=1.21e-06 nrd=0.578824 nrs=0.211765 sa=1.94353e-06 sb=4.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.8e-14 panw10=0 $X=136170 $Y=45240 $D=111
M8410 78 112 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.16e-13 pd=1.66e-06 ps=3.24e-06 nrd=0.138462 nrs=0.246154 sa=3.2e-07 sb=1.66215e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=33210 $Y=35510 $D=111
M8411 VDD 112 78 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=2.34e-13 pd=1.66e-06 ps=1.66e-06 nrd=0.138462 nrs=0.138462 sa=8e-07 sb=1.18215e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=33690 $Y=35510 $D=111
M8412 78 112 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.45898e-13 as=2.34e-13 pd=1.82881e-06 ps=1.66e-06 nrd=0.145502 nrs=0.138462 sa=1.28e-06 sb=7.02154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=34170 $Y=35510 $D=111
M8413 VDD 112 78 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=2.00502e-13 pd=2.76e-06 ps=1.49119e-06 nrd=0.301887 nrs=0.178446 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=34650 $Y=35510 $D=111
M8414 123 112 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.16e-13 pd=1.66e-06 ps=3.24e-06 nrd=0.138462 nrs=0.246154 sa=3.2e-07 sb=1.66215e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=34410 $Y=42710 $D=111
M8415 VDD 112 123 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=2.34e-13 pd=1.66e-06 ps=1.66e-06 nrd=0.138462 nrs=0.138462 sa=8e-07 sb=1.18215e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=34890 $Y=42710 $D=111
M8416 123 112 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.45898e-13 as=2.34e-13 pd=1.82881e-06 ps=1.66e-06 nrd=0.145502 nrs=0.138462 sa=1.28e-06 sb=7.02154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=35370 $Y=42710 $D=111
M8417 VDD 112 123 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=2.00502e-13 pd=2.76e-06 ps=1.49119e-06 nrd=0.301887 nrs=0.178446 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=35850 $Y=42710 $D=111
M8418 278 236 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.16e-13 pd=1.66e-06 ps=3.24e-06 nrd=0.138462 nrs=0.246154 sa=3.2e-07 sb=1.66215e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=58410 $Y=30390 $D=111
M8419 VDD 236 278 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=2.34e-13 pd=1.66e-06 ps=1.66e-06 nrd=0.138462 nrs=0.138462 sa=8e-07 sb=1.18215e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=58890 $Y=30390 $D=111
M8420 278 236 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.45898e-13 as=2.34e-13 pd=1.82881e-06 ps=1.66e-06 nrd=0.145502 nrs=0.138462 sa=1.28e-06 sb=7.02154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=59370 $Y=30390 $D=111
M8421 VDD 236 278 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=2.00502e-13 pd=2.76e-06 ps=1.49119e-06 nrd=0.301887 nrs=0.178446 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=59850 $Y=30630 $D=111
M8422 231 263 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.16e-13 pd=1.66e-06 ps=3.24e-06 nrd=0.138462 nrs=0.246154 sa=3.2e-07 sb=1.66215e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=61210 $Y=30390 $D=111
M8423 VDD 263 231 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=2.34e-13 pd=1.66e-06 ps=1.66e-06 nrd=0.138462 nrs=0.138462 sa=8e-07 sb=1.18215e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=61690 $Y=30390 $D=111
M8424 231 263 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.45898e-13 as=2.34e-13 pd=1.82881e-06 ps=1.66e-06 nrd=0.145502 nrs=0.138462 sa=1.28e-06 sb=7.02154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=62170 $Y=30390 $D=111
M8425 VDD 263 231 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=2.00502e-13 pd=2.76e-06 ps=1.49119e-06 nrd=0.301887 nrs=0.178446 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=62650 $Y=30630 $D=111
M8426 301 284 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.16e-13 pd=1.66e-06 ps=3.24e-06 nrd=0.138462 nrs=0.246154 sa=3.2e-07 sb=1.66215e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=75610 $Y=37590 $D=111
M8427 VDD 284 301 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=2.34e-13 pd=1.66e-06 ps=1.66e-06 nrd=0.138462 nrs=0.138462 sa=8e-07 sb=1.18215e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=76090 $Y=37590 $D=111
M8428 301 284 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.45898e-13 as=2.34e-13 pd=1.82881e-06 ps=1.66e-06 nrd=0.145502 nrs=0.138462 sa=1.28e-06 sb=7.02154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=76570 $Y=37590 $D=111
M8429 VDD 284 301 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=2.00502e-13 pd=2.76e-06 ps=1.49119e-06 nrd=0.301887 nrs=0.178446 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=77050 $Y=37830 $D=111
M8430 523 503 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=4.16e-13 pd=1.66e-06 ps=3.24e-06 nrd=0.138462 nrs=0.246154 sa=3.2e-07 sb=1.66215e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=131210 $Y=64310 $D=111
M8431 VDD 503 523 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.34e-13 as=2.34e-13 pd=1.66e-06 ps=1.66e-06 nrd=0.138462 nrs=0.138462 sa=8e-07 sb=1.18215e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=131690 $Y=64310 $D=111
M8432 523 503 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.45898e-13 as=2.34e-13 pd=1.82881e-06 ps=1.66e-06 nrd=0.145502 nrs=0.138462 sa=1.28e-06 sb=7.02154e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=132170 $Y=64310 $D=111
M8433 VDD 503 523 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=2.00502e-13 pd=2.76e-06 ps=1.49119e-06 nrd=0.301887 nrs=0.178446 sa=1.76e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=132650 $Y=64310 $D=111
M8434 3773 49 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=18430 $Y=28310 $D=111
M8435 VDD 49 3773 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=18910 $Y=28310 $D=111
M8436 3772 3773 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=19350 $Y=28310 $D=111
M8437 VDD 3773 3772 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=19830 $Y=28310 $D=111
M8438 3771 78 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=20270 $Y=28310 $D=111
M8439 3772 3771 57 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=21230 $Y=28510 $D=111
M8440 57 3771 3772 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=21710 $Y=28510 $D=111
M8441 3773 78 57 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=22190 $Y=28530 $D=111
M8442 57 78 3773 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=22670 $Y=28530 $D=111
M8443 3776 127 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=25630 $Y=35510 $D=111
M8444 VDD 127 3776 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=26110 $Y=35510 $D=111
M8445 3775 3776 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=26550 $Y=35510 $D=111
M8446 VDD 3776 3775 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=27030 $Y=35510 $D=111
M8447 3774 123 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=27470 $Y=35510 $D=111
M8448 3775 3774 107 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=28430 $Y=35710 $D=111
M8449 107 3774 3775 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=28910 $Y=35710 $D=111
M8450 3776 123 107 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=29390 $Y=35730 $D=111
M8451 107 123 3776 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=29870 $Y=35730 $D=111
M8452 3779 136 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=32030 $Y=45310 $D=111
M8453 VDD 136 3779 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=32510 $Y=45310 $D=111
M8454 3778 3779 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=32950 $Y=45310 $D=111
M8455 VDD 3779 3778 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=33430 $Y=45310 $D=111
M8456 3777 123 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=33870 $Y=45470 $D=111
M8457 3778 3777 131 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=34830 $Y=45110 $D=111
M8458 131 3777 3778 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=35310 $Y=45110 $D=111
M8459 3779 123 131 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=35790 $Y=45090 $D=111
M8460 131 123 3779 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=36270 $Y=45090 $D=111
M8461 3782 141 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=34030 $Y=30910 $D=111
M8462 VDD 141 3782 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=34510 $Y=30910 $D=111
M8463 3781 3782 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=34950 $Y=30910 $D=111
M8464 VDD 3782 3781 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=35430 $Y=30910 $D=111
M8465 3780 78 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=35870 $Y=31070 $D=111
M8466 3781 3780 142 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=36830 $Y=30710 $D=111
M8467 142 3780 3781 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=37310 $Y=30710 $D=111
M8468 3782 78 142 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=37790 $Y=30690 $D=111
M8469 142 78 3782 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=38270 $Y=30690 $D=111
M8470 3785 127 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=36030 $Y=35510 $D=111
M8471 VDD 127 3785 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=36510 $Y=35510 $D=111
M8472 3784 3785 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=36950 $Y=35510 $D=111
M8473 VDD 3785 3784 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=37430 $Y=35510 $D=111
M8474 3783 123 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=37870 $Y=35510 $D=111
M8475 3784 3783 893 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=38830 $Y=35710 $D=111
M8476 893 3783 3784 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=39310 $Y=35710 $D=111
M8477 3785 123 893 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=39790 $Y=35730 $D=111
M8478 893 123 3785 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=40270 $Y=35730 $D=111
M8479 3788 157 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=40030 $Y=42710 $D=111
M8480 VDD 157 3788 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=40510 $Y=42710 $D=111
M8481 3787 3788 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=40950 $Y=42710 $D=111
M8482 VDD 3788 3787 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=41430 $Y=42710 $D=111
M8483 3786 163 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=41870 $Y=42710 $D=111
M8484 3787 3786 166 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=42830 $Y=42910 $D=111
M8485 166 3786 3787 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=43310 $Y=42910 $D=111
M8486 3788 163 166 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=43790 $Y=42930 $D=111
M8487 166 163 3788 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=44270 $Y=42930 $D=111
M8488 3791 157 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=40430 $Y=52510 $D=111
M8489 VDD 157 3791 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=40910 $Y=52510 $D=111
M8490 3790 3791 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=41350 $Y=52510 $D=111
M8491 VDD 3791 3790 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=41830 $Y=52510 $D=111
M8492 3789 78 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=42270 $Y=52670 $D=111
M8493 3790 3789 174 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=43230 $Y=52310 $D=111
M8494 174 3789 3790 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=43710 $Y=52310 $D=111
M8495 3791 78 174 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=44190 $Y=52290 $D=111
M8496 174 78 3791 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=44670 $Y=52290 $D=111
M8497 3794 78 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=43630 $Y=57110 $D=111
M8498 VDD 78 3794 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=44110 $Y=57110 $D=111
M8499 3793 3794 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=44550 $Y=57110 $D=111
M8500 VDD 3794 3793 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=45030 $Y=57110 $D=111
M8501 3792 186 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=45470 $Y=57110 $D=111
M8502 3793 3792 181 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=46430 $Y=57310 $D=111
M8503 181 3792 3793 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=46910 $Y=57310 $D=111
M8504 3794 186 181 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=47390 $Y=57330 $D=111
M8505 181 186 3794 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=47870 $Y=57330 $D=111
M8506 3797 171 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=45630 $Y=52510 $D=111
M8507 VDD 171 3797 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=46110 $Y=52510 $D=111
M8508 3796 3797 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=46550 $Y=52510 $D=111
M8509 VDD 3797 3796 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=47030 $Y=52510 $D=111
M8510 3795 78 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=47470 $Y=52670 $D=111
M8511 3796 3795 179 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=48430 $Y=52310 $D=111
M8512 179 3795 3796 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=48910 $Y=52310 $D=111
M8513 3797 78 179 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=49390 $Y=52290 $D=111
M8514 179 78 3797 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=49870 $Y=52290 $D=111
M8515 3800 240 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=74830 $Y=28310 $D=111
M8516 VDD 240 3800 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=75310 $Y=28310 $D=111
M8517 3799 3800 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=75750 $Y=28310 $D=111
M8518 VDD 3800 3799 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=76230 $Y=28310 $D=111
M8519 3798 287 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=76670 $Y=28310 $D=111
M8520 3799 3798 280 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=77630 $Y=28510 $D=111
M8521 280 3798 3799 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=78110 $Y=28510 $D=111
M8522 3800 287 280 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=78590 $Y=28530 $D=111
M8523 280 287 3800 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=79070 $Y=28530 $D=111
M8524 3803 240 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=74830 $Y=30910 $D=111
M8525 VDD 240 3803 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=75310 $Y=30910 $D=111
M8526 3802 3803 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=75750 $Y=30910 $D=111
M8527 VDD 3803 3802 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=76230 $Y=30910 $D=111
M8528 3801 254 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=76670 $Y=31070 $D=111
M8529 3802 3801 293 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=77630 $Y=30710 $D=111
M8530 293 3801 3802 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=78110 $Y=30710 $D=111
M8531 3803 254 293 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=78590 $Y=30690 $D=111
M8532 293 254 3803 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=79070 $Y=30690 $D=111
M8533 3806 157 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=79230 $Y=45310 $D=111
M8534 VDD 157 3806 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=79710 $Y=45310 $D=111
M8535 3805 3806 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=80150 $Y=45310 $D=111
M8536 VDD 3806 3805 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=80630 $Y=45310 $D=111
M8537 3804 307 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=81070 $Y=45470 $D=111
M8538 3805 3804 319 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=82030 $Y=45110 $D=111
M8539 319 3804 3805 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=82510 $Y=45110 $D=111
M8540 3806 307 319 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=82990 $Y=45090 $D=111
M8541 319 307 3806 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=83470 $Y=45090 $D=111
M8542 3809 186 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=80430 $Y=57110 $D=111
M8543 VDD 186 3809 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=80910 $Y=57110 $D=111
M8544 3808 3809 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=81350 $Y=57110 $D=111
M8545 VDD 3809 3808 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=81830 $Y=57110 $D=111
M8546 3807 307 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=82270 $Y=57110 $D=111
M8547 3808 3807 314 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=83230 $Y=57310 $D=111
M8548 314 3807 3808 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=83710 $Y=57310 $D=111
M8549 3809 307 314 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=84190 $Y=57330 $D=111
M8550 314 307 3809 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=84670 $Y=57330 $D=111
M8551 3812 354 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=84030 $Y=35510 $D=111
M8552 VDD 354 3812 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=84510 $Y=35510 $D=111
M8553 3811 3812 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=84950 $Y=35510 $D=111
M8554 VDD 3812 3811 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=85430 $Y=35510 $D=111
M8555 3810 192 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=85870 $Y=35510 $D=111
M8556 3811 3810 328 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=86830 $Y=35710 $D=111
M8557 328 3810 3811 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=87310 $Y=35710 $D=111
M8558 3812 192 328 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=87790 $Y=35730 $D=111
M8559 328 192 3812 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=88270 $Y=35730 $D=111
M8560 3815 171 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=84430 $Y=45310 $D=111
M8561 VDD 171 3815 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=84910 $Y=45310 $D=111
M8562 3814 3815 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=85350 $Y=45310 $D=111
M8563 VDD 3815 3814 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=85830 $Y=45310 $D=111
M8564 3813 307 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=86270 $Y=45470 $D=111
M8565 3814 3813 327 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=87230 $Y=45110 $D=111
M8566 327 3813 3814 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=87710 $Y=45110 $D=111
M8567 3815 307 327 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=88190 $Y=45090 $D=111
M8568 327 307 3815 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=88670 $Y=45090 $D=111
M8569 3818 176 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=88430 $Y=38110 $D=111
M8570 VDD 176 3818 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=88910 $Y=38110 $D=111
M8571 3817 3818 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=89350 $Y=38110 $D=111
M8572 VDD 3818 3817 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=89830 $Y=38110 $D=111
M8573 3816 354 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=90270 $Y=38270 $D=111
M8574 3817 3816 343 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=91230 $Y=37910 $D=111
M8575 343 3816 3817 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=91710 $Y=37910 $D=111
M8576 3818 354 343 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=92190 $Y=37890 $D=111
M8577 343 354 3818 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=92670 $Y=37890 $D=111
M8578 3821 538 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=104830 $Y=49910 $D=111
M8579 VDD 538 3821 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=105310 $Y=49910 $D=111
M8580 3820 3821 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=105750 $Y=49910 $D=111
M8581 VDD 3821 3820 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=106230 $Y=49910 $D=111
M8582 3819 395 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=106670 $Y=49910 $D=111
M8583 3820 3819 406 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=107630 $Y=50110 $D=111
M8584 406 3819 3820 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=108110 $Y=50110 $D=111
M8585 3821 395 406 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=108590 $Y=50130 $D=111
M8586 406 395 3821 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=109070 $Y=50130 $D=111
M8587 3824 520 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.652e-13 pd=1.14e-06 ps=2.24e-06 nrd=0.230769 nrs=0.435897 sa=3.4e-07 sb=1.92615e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=127630 $Y=52510 $D=111
M8588 VDD 520 3824 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.80757e-13 as=1.404e-13 pd=1.70413e-06 ps=1.14e-06 nrd=0.297101 nrs=0.230769 sa=8.2e-07 sb=1.57333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=128110 $Y=52510 $D=111
M8589 3823 3824 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.80757e-13 pd=1.14e-06 ps=1.70413e-06 nrd=0.230769 nrs=0.297101 sa=1.26e-06 sb=1.13333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=128550 $Y=52510 $D=111
M8590 VDD 3824 3823 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.00386e-13 as=1.404e-13 pd=1.86643e-06 ps=1.14e-06 nrd=0.329365 nrs=0.230769 sa=1.74e-06 sb=6.53333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=129030 $Y=52510 $D=111
M8591 3822 545 VDD VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.984e-13 as=1.59281e-13 pd=1.88e-06 ps=1.48357e-06 nrd=0.516129 nrs=0.414363 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.44e-14 panw9=0 panw10=0 $X=129470 $Y=52670 $D=111
M8592 3823 3822 466 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.496e-13 pd=1.14e-06 ps=2.2e-06 nrd=0.230769 nrs=0.410256 sa=3.2e-07 sb=1.73282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=130430 $Y=52310 $D=111
M8593 466 3822 3823 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.414e-13 as=1.404e-13 pd=1.16e-06 ps=1.14e-06 nrd=0.232413 nrs=0.230769 sa=8e-07 sb=1.25282e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=130910 $Y=52310 $D=111
M8594 3824 545 466 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=1.414e-13 pd=1.14e-06 ps=1.16e-06 nrd=0.230769 nrs=0.232413 sa=1.25333e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=131390 $Y=52290 $D=111
M8595 466 545 3824 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=1.404e-13 pd=2.2e-06 ps=1.14e-06 nrd=0.410256 nrs=0.230769 sa=1.73333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=9.6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=131870 $Y=52290 $D=111
M8596 30 21 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=12400 $Y=37590 $D=111
M8597 VDD 17 30 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=12880 $Y=37590 $D=111
M8598 30 17 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=13360 $Y=37590 $D=111
M8599 VDD 21 30 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=13840 $Y=37590 $D=111
M8600 59 48 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=12800 $Y=51990 $D=111
M8601 VDD 14 59 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=13280 $Y=51990 $D=111
M8602 59 14 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=13760 $Y=51990 $D=111
M8603 VDD 48 59 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=14240 $Y=51990 $D=111
M8604 53 800 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=14800 $Y=35520 $D=111
M8605 VDD 34 53 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=15280 $Y=35520 $D=111
M8606 53 34 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=15760 $Y=35520 $D=111
M8607 VDD 800 53 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=16240 $Y=35520 $D=111
M8608 98 96 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=27200 $Y=59190 $D=111
M8609 VDD 73 98 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=27680 $Y=59190 $D=111
M8610 98 73 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=28160 $Y=59190 $D=111
M8611 VDD 96 98 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=28640 $Y=59190 $D=111
M8612 168 163 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=38800 $Y=21120 $D=111
M8613 VDD 148 168 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=39280 $Y=21120 $D=111
M8614 168 148 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=39760 $Y=21120 $D=111
M8615 VDD 163 168 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=40240 $Y=21120 $D=111
M8616 182 163 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=43200 $Y=23190 $D=111
M8617 VDD 148 182 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=43680 $Y=23190 $D=111
M8618 182 148 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=44160 $Y=23190 $D=111
M8619 VDD 163 182 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=44640 $Y=23190 $D=111
M8620 169 177 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=48400 $Y=15990 $D=111
M8621 VDD 143 169 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=48880 $Y=15990 $D=111
M8622 169 143 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=49360 $Y=15990 $D=111
M8623 VDD 177 169 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=49840 $Y=15990 $D=111
M8624 242 285 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=64800 $Y=30390 $D=111
M8625 VDD 278 242 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=65280 $Y=30390 $D=111
M8626 242 278 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=65760 $Y=30390 $D=111
M8627 VDD 285 242 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=66240 $Y=30390 $D=111
M8628 246 245 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=65600 $Y=49920 $D=111
M8629 VDD 213 246 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=66080 $Y=49920 $D=111
M8630 246 213 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=66560 $Y=49920 $D=111
M8631 VDD 245 246 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=67040 $Y=49920 $D=111
M8632 282 291 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=73600 $Y=35520 $D=111
M8633 VDD 278 282 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=74080 $Y=35520 $D=111
M8634 282 278 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=74560 $Y=35520 $D=111
M8635 VDD 291 282 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=75040 $Y=35520 $D=111
M8636 358 347 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=79600 $Y=73590 $D=111
M8637 VDD 308 358 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=80080 $Y=73590 $D=111
M8638 358 308 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=80560 $Y=73590 $D=111
M8639 VDD 347 358 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=81040 $Y=73590 $D=111
M8640 330 278 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=80400 $Y=37590 $D=111
M8641 VDD 301 330 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=80880 $Y=37590 $D=111
M8642 330 301 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=81360 $Y=37590 $D=111
M8643 VDD 278 330 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=81840 $Y=37590 $D=111
M8644 476 401 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=106000 $Y=64320 $D=111
M8645 VDD 392 476 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=106480 $Y=64320 $D=111
M8646 476 392 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=106960 $Y=64320 $D=111
M8647 VDD 401 476 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=107440 $Y=64320 $D=111
M8648 405 836 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=115200 $Y=30390 $D=111
M8649 VDD 427 405 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=115680 $Y=30390 $D=111
M8650 405 427 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=116160 $Y=30390 $D=111
M8651 VDD 836 405 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=116640 $Y=30390 $D=111
M8652 496 473 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=6.49359e-13 pd=1.65e-06 ps=2.73315e-06 nrd=0.139535 nrs=0.390216 sa=7.6e-07 sb=1.76e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=128000 $Y=73590 $D=111
M8653 VDD 490 496 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.24e-06 sb=1.28e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=128480 $Y=73590 $D=111
M8654 496 490 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.322e-13 pd=1.65e-06 ps=1.65e-06 nrd=0.139535 nrs=0.139535 sa=1.72e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=128960 $Y=73590 $D=111
M8655 VDD 473 496 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=129440 $Y=73590 $D=111
M8656 284 216 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=57230 $Y=42710 $D=111
M8657 VDD 206 284 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=57710 $Y=42710 $D=111
M8658 284 206 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=58190 $Y=42710 $D=111
M8659 VDD 216 284 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.76e-06 sb=1.54e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=58670 $Y=42710 $D=111
M8660 284 216 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.304e-13 pd=1.72e-06 ps=1.64e-06 nrd=0.171875 nrs=0.140625 sa=2e-06 sb=1.06e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=59150 $Y=42710 $D=111
M8661 VDD 206 284 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.07867e-13 as=2.816e-13 pd=2.76e-06 ps=1.72e-06 nrd=0.309977 nrs=0.171875 sa=2e-06 sb=5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=59710 $Y=42710 $D=111
M8662 232 278 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=80030 $Y=35510 $D=111
M8663 VDD 304 232 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=80510 $Y=35510 $D=111
M8664 232 304 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=80990 $Y=35510 $D=111
M8665 VDD 278 232 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.76e-06 sb=1.54e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=81470 $Y=35510 $D=111
M8666 232 278 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.304e-13 pd=1.72e-06 ps=1.64e-06 nrd=0.171875 nrs=0.140625 sa=2e-06 sb=1.06e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=81950 $Y=35510 $D=111
M8667 VDD 304 232 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.07867e-13 as=2.816e-13 pd=2.76e-06 ps=1.72e-06 nrd=0.309977 nrs=0.171875 sa=2e-06 sb=5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=82510 $Y=35510 $D=111
M8668 846 460 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=126430 $Y=64310 $D=111
M8669 VDD 443 846 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=126910 $Y=64310 $D=111
M8670 846 443 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.28e-06 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=127390 $Y=64310 $D=111
M8671 VDD 460 846 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.76e-06 sb=1.54e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=127870 $Y=64310 $D=111
M8672 846 460 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.816e-13 as=2.304e-13 pd=1.72e-06 ps=1.64e-06 nrd=0.171875 nrs=0.140625 sa=2e-06 sb=1.06e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=128350 $Y=64310 $D=111
M8673 VDD 443 846 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.07867e-13 as=2.816e-13 pd=2.76e-06 ps=1.72e-06 nrd=0.309977 nrs=0.171875 sa=2e-06 sb=5e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=128910 $Y=64310 $D=111
M8674 VDD 228 3882 VDD lppfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.19429e-13 as=3.84e-13 pd=1.67143e-06 ps=3.04e-06 nrd=0.152381 nrs=0.266667 sa=3.2e-07 sb=1.65533e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=56920 $Y=57110 $D=111
M8675 3883 218 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.04e-13 as=1.90171e-13 pd=1.24e-06 ps=1.44857e-06 nrd=0.0961538 nrs=0.175824 sa=8e-07 sb=1.81154e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=57400 $Y=57110 $D=111
M8676 211 3882 3883 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.005e-13 as=1.04e-13 pd=1.54e-06 ps=1.24e-06 nrd=0.185374 nrs=0.0961538 sa=1.12e-06 sb=1.69923e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=57720 $Y=57110 $D=111
M8677 3884 3882 211 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.04e-13 as=2.005e-13 pd=1.24e-06 ps=1.54e-06 nrd=0.0961538 nrs=0.185374 sa=1.42096e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=58200 $Y=57250 $D=111
M8678 VDD 218 3884 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.04e-13 pd=1.4e-06 ps=1.24e-06 nrd=0.173077 nrs=0.0961538 sa=1.74096e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=58520 $Y=57250 $D=111
M8679 3885 218 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.04e-13 as=1.872e-13 pd=1.24e-06 ps=1.4e-06 nrd=0.0961538 nrs=0.173077 sa=1.87481e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=59000 $Y=57250 $D=111
M8680 211 3882 3885 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.04e-13 pd=2.72e-06 ps=1.24e-06 nrd=0.307692 nrs=0.0961538 sa=1.91788e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=59320 $Y=57250 $D=111
M8681 VDD 466 3886 VDD lppfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.19429e-13 as=3.84e-13 pd=1.67143e-06 ps=3.04e-06 nrd=0.152381 nrs=0.266667 sa=3.2e-07 sb=1.65533e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=124120 $Y=52090 $D=111
M8682 3887 485 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.04e-13 as=1.90171e-13 pd=1.24e-06 ps=1.44857e-06 nrd=0.0961538 nrs=0.175824 sa=8e-07 sb=1.81154e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=124600 $Y=52250 $D=111
M8683 475 3886 3887 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.005e-13 as=1.04e-13 pd=1.54e-06 ps=1.24e-06 nrd=0.185374 nrs=0.0961538 sa=1.12e-06 sb=1.69923e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=124920 $Y=52250 $D=111
M8684 3888 3886 475 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.04e-13 as=2.005e-13 pd=1.24e-06 ps=1.54e-06 nrd=0.0961538 nrs=0.185374 sa=1.42096e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=125400 $Y=52110 $D=111
M8685 VDD 485 3888 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.872e-13 as=1.04e-13 pd=1.4e-06 ps=1.24e-06 nrd=0.173077 nrs=0.0961538 sa=1.74096e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=125720 $Y=52110 $D=111
M8686 3889 485 VDD VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.04e-13 as=1.872e-13 pd=1.24e-06 ps=1.4e-06 nrd=0.0961538 nrs=0.173077 sa=1.87481e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=126200 $Y=52110 $D=111
M8687 475 3886 3889 VDD lppfet w=1.04e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.328e-13 as=1.04e-13 pd=2.72e-06 ps=1.24e-06 nrd=0.307692 nrs=0.0961538 sa=1.91788e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=126520 $Y=52110 $D=111
M8688 3891 8 3890 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3e-13 as=4.16e-13 pd=1.5e-06 ps=3.24e-06 nrd=0.0769231 nrs=0.246154 sa=3.2e-07 sb=1.624e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.02e-13 panw9=1.26e-13 panw10=2.4e-14 $X=9000 $Y=37590 $D=111
M8689 VDD 17 3891 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.92319e-13 as=1.3e-13 pd=1.81458e-06 ps=1.5e-06 nrd=0.17297 nrs=0.0769231 sa=6.4e-07 sb=1.304e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-13 panw10=2.4e-14 $X=9320 $Y=37590 $D=111
M8690 14 3890 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.41398e-13 as=2.92319e-13 pd=1.75447e-06 ps=1.81458e-06 nrd=0.142839 nrs=0.17297 sa=1.2e-06 sb=7.44e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.8e-13 $X=9880 $Y=37590 $D=111
M8691 VDD 3890 14 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.712e-13 as=2.15402e-13 pd=2.96e-06 ps=1.56553e-06 nrd=0.275862 nrs=0.160078 sa=1.68e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=10360 $Y=37730 $D=111
M8692 3893 156 3892 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3e-13 as=4.16e-13 pd=1.5e-06 ps=3.24e-06 nrd=0.0769231 nrs=0.246154 sa=3.2e-07 sb=1.624e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=36600 $Y=51990 $D=111
M8693 VDD 146 3893 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.92319e-13 as=1.3e-13 pd=1.81458e-06 ps=1.5e-06 nrd=0.17297 nrs=0.0769231 sa=6.4e-07 sb=1.304e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=36920 $Y=51990 $D=111
M8694 138 3892 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.41398e-13 as=2.92319e-13 pd=1.75447e-06 ps=1.81458e-06 nrd=0.142839 nrs=0.17297 sa=1.2e-06 sb=7.44e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=37480 $Y=51990 $D=111
M8695 VDD 3892 138 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.712e-13 as=2.15402e-13 pd=2.96e-06 ps=1.56553e-06 nrd=0.275862 nrs=0.160078 sa=1.68e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=37960 $Y=52130 $D=111
M8696 3895 146 3894 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3e-13 as=4.16e-13 pd=1.5e-06 ps=3.24e-06 nrd=0.0769231 nrs=0.246154 sa=3.2e-07 sb=1.624e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=39800 $Y=57110 $D=111
M8697 VDD 156 3895 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.92319e-13 as=1.3e-13 pd=1.81458e-06 ps=1.5e-06 nrd=0.17297 nrs=0.0769231 sa=6.4e-07 sb=1.304e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=40120 $Y=57110 $D=111
M8698 160 3894 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.41398e-13 as=2.92319e-13 pd=1.75447e-06 ps=1.81458e-06 nrd=0.142839 nrs=0.17297 sa=1.2e-06 sb=7.44e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=40680 $Y=57110 $D=111
M8699 VDD 3894 160 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.712e-13 as=2.15402e-13 pd=2.96e-06 ps=1.56553e-06 nrd=0.275862 nrs=0.160078 sa=1.68e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=41160 $Y=57110 $D=111
M8700 3897 248 3896 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3e-13 as=4.16e-13 pd=1.5e-06 ps=3.24e-06 nrd=0.0769231 nrs=0.246154 sa=3.2e-07 sb=1.624e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=75800 $Y=57110 $D=111
M8701 VDD 239 3897 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.92319e-13 as=1.3e-13 pd=1.81458e-06 ps=1.5e-06 nrd=0.17297 nrs=0.0769231 sa=6.4e-07 sb=1.304e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=76120 $Y=57110 $D=111
M8702 315 3896 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.41398e-13 as=2.92319e-13 pd=1.75447e-06 ps=1.81458e-06 nrd=0.142839 nrs=0.17297 sa=1.2e-06 sb=7.44e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=76680 $Y=57110 $D=111
M8703 VDD 3896 315 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.712e-13 as=2.15402e-13 pd=2.96e-06 ps=1.56553e-06 nrd=0.275862 nrs=0.160078 sa=1.68e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=77160 $Y=57110 $D=111
M8704 3899 463 3898 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3e-13 as=4.16e-13 pd=1.5e-06 ps=3.24e-06 nrd=0.0769231 nrs=0.246154 sa=3.2e-07 sb=1.624e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=121400 $Y=51990 $D=111
M8705 VDD 457 3899 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.92319e-13 as=1.3e-13 pd=1.81458e-06 ps=1.5e-06 nrd=0.17297 nrs=0.0769231 sa=6.4e-07 sb=1.304e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=121720 $Y=51990 $D=111
M8706 460 3898 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.41398e-13 as=2.92319e-13 pd=1.75447e-06 ps=1.81458e-06 nrd=0.142839 nrs=0.17297 sa=1.2e-06 sb=7.44e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=122280 $Y=51990 $D=111
M8707 VDD 3898 460 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.712e-13 as=2.15402e-13 pd=2.96e-06 ps=1.56553e-06 nrd=0.275862 nrs=0.160078 sa=1.68e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=122760 $Y=52130 $D=111
M8708 799 40 VDD VDD lppfet w=9.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.71e-13 as=3.04e-13 pd=1.31e-06 ps=2.54e-06 nrd=0.189474 nrs=0.336842 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3e-14 panw10=0 $X=14090 $Y=21110 $D=111
M8709 VDD 40 799 VDD lppfet w=9.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.23e-13 as=1.71e-13 pd=2.58e-06 ps=1.31e-06 nrd=0.357895 nrs=0.189474 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3e-14 panw10=0 $X=14570 $Y=21110 $D=111
M8710 177 188 VDD VDD lppfet w=9.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.71e-13 as=3.04e-13 pd=1.31e-06 ps=2.54e-06 nrd=0.189474 nrs=0.336842 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3e-14 panw10=0 $X=46090 $Y=16340 $D=111
M8711 VDD 188 177 VDD lppfet w=9.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.23e-13 as=1.71e-13 pd=2.58e-06 ps=1.31e-06 nrd=0.357895 nrs=0.189474 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3e-14 panw10=0 $X=46570 $Y=16340 $D=111
M8712 377 368 VDD VDD lppfet w=9.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.71e-13 as=3.04e-13 pd=1.31e-06 ps=2.54e-06 nrd=0.189474 nrs=0.336842 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3e-14 panw10=0 $X=94490 $Y=16340 $D=111
M8713 VDD 368 377 VDD lppfet w=9.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.23e-13 as=1.71e-13 pd=2.58e-06 ps=1.31e-06 nrd=0.357895 nrs=0.189474 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3e-14 panw10=0 $X=94970 $Y=16340 $D=111
M8714 836 441 VDD VDD lppfet w=9.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.71e-13 as=3.04e-13 pd=1.31e-06 ps=2.54e-06 nrd=0.189474 nrs=0.336842 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3e-14 panw10=0 $X=112890 $Y=30740 $D=111
M8715 VDD 441 836 VDD lppfet w=9.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.23e-13 as=1.71e-13 pd=2.58e-06 ps=1.31e-06 nrd=0.357895 nrs=0.189474 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3e-14 panw10=0 $X=113370 $Y=30740 $D=111
M8716 467 432 VDD VDD lppfet w=9.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.71e-13 as=3.04e-13 pd=1.31e-06 ps=2.54e-06 nrd=0.189474 nrs=0.336842 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3e-14 panw10=0 $X=119290 $Y=59540 $D=111
M8717 VDD 432 467 VDD lppfet w=9.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.23e-13 as=1.71e-13 pd=2.58e-06 ps=1.31e-06 nrd=0.357895 nrs=0.189474 sa=8e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3e-14 panw10=0 $X=119770 $Y=59540 $D=111
M8718 VDD 910 3902 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.41899e-13 as=4.096e-13 pd=2.10211e-06 ps=3.2e-06 nrd=0.147644 nrs=0.25 sa=3.2e-07 sb=1.15758e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=110410 $Y=44790 $D=111
M8719 3900 3902 VDD VDD lppfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.6959e-13 as=1.70085e-13 pd=1.36627e-06 ps=1.47805e-06 nrd=0.209371 nrs=0.209982 sa=7.47556e-07 sb=1.26889e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=110850 $Y=45190 $D=111
M8720 3906 3901 3900 VDD lppfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.03873e-13 as=1.4321e-13 pd=1.54413e-06 ps=1.15373e-06 nrd=0.352966 nrs=0.247939 sa=1.22526e-06 sb=9.71053e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=7.2e-15 panw10=0 $X=111330 $Y=45330 $D=111
M8721 3901 3900 3906 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.1191e-13 as=1.34127e-13 pd=9.21348e-07 ps=1.01587e-06 nrd=0.44764 nrs=0.536508 sa=1.8576e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=111970 $Y=45590 $D=111
M8722 VDD 436 3901 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.39692e-13 as=2.8649e-13 pd=3.16718e-06 ps=2.35865e-06 nrd=0.207332 nrs=0.17486 sa=9.4875e-07 sb=2.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=112450 $Y=44810 $D=111
M8723 3904 3902 3901 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.00317e-13 as=1.6e-13 pd=8.88889e-07 ps=1.64e-06 nrd=0.40127 nrs=0.64 sa=3.2e-07 sb=8.344e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=8.4e-15 panw9=0 panw10=0 $X=113270 $Y=45470 $D=111
M8724 3902 3901 3904 VDD lppfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.77816e-13 as=1.52483e-13 pd=1.60444e-06 ps=1.35111e-06 nrd=0.307853 nrs=0.263993 sa=6.22105e-07 sb=9.05789e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=113750 $Y=45210 $D=111
M8725 3905 3904 3902 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9e-14 as=1.16984e-13 pd=8.6e-07 ps=1.05556e-06 nrd=0.36 nrs=0.467937 sa=5.896e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=4.08e-14 panw10=0 $X=114230 $Y=45000 $D=111
M8726 3903 3906 3905 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.5e-13 as=9e-14 pd=1.1e-06 ps=8.6e-07 nrd=0.6 nrs=0.36 sa=1.0696e-06 sb=9.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=4.08e-14 panw10=0 $X=114710 $Y=45000 $D=111
M8727 VDD 451 3903 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.6e-13 as=1.5e-13 pd=1.71795e-06 ps=1.1e-06 nrd=0.64 nrs=0.6 sa=1.7608e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=4.08e-14 panw10=0 $X=115430 $Y=45000 $D=111
M8728 3907 3903 3904 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9e-14 as=1.6e-13 pd=8.6e-07 ps=1.64e-06 nrd=0.36 nrs=0.64 sa=3.2e-07 sb=7.856e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=116390 $Y=45260 $D=111
M8729 3906 451 3907 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.528e-13 as=9e-14 pd=1.64e-06 ps=8.6e-07 nrd=0.6112 nrs=0.36 sa=8e-07 sb=3.056e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=116870 $Y=45260 $D=111
M8730 VDD 3905 480 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=3.092e-13 pd=1.64e-06 ps=3.42e-06 nrd=0.140625 nrs=0.188721 sa=2.2625e-07 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=117690 $Y=44810 $D=111
M8731 457 3907 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=7.0625e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=118170 $Y=44810 $D=111
M8732 VDD 839 3910 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.41899e-13 as=4.096e-13 pd=2.10211e-06 ps=3.2e-06 nrd=0.147644 nrs=0.25 sa=3.2e-07 sb=1.15758e-06 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=118410 $Y=42730 $D=111
M8733 3908 3910 VDD VDD lppfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.6959e-13 as=1.70085e-13 pd=1.36627e-06 ps=1.47805e-06 nrd=0.209371 nrs=0.209982 sa=7.47556e-07 sb=1.26889e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=118850 $Y=42710 $D=111
M8734 3914 3909 3908 VDD lppfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.03873e-13 as=1.4321e-13 pd=1.54413e-06 ps=1.15373e-06 nrd=0.352966 nrs=0.247939 sa=1.22526e-06 sb=9.71053e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=7.2e-15 panw10=0 $X=119330 $Y=42710 $D=111
M8735 3909 3908 3914 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.1191e-13 as=1.34127e-13 pd=9.21348e-07 ps=1.01587e-06 nrd=0.44764 nrs=0.536508 sa=1.8576e-06 sb=6.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=119970 $Y=42710 $D=111
M8736 VDD 444 3909 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.39692e-13 as=2.8649e-13 pd=3.16718e-06 ps=2.35865e-06 nrd=0.207332 nrs=0.17486 sa=9.4875e-07 sb=2.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=120450 $Y=42710 $D=111
M8737 3912 3910 3909 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.00317e-13 as=1.6e-13 pd=8.88889e-07 ps=1.64e-06 nrd=0.40127 nrs=0.64 sa=3.2e-07 sb=8.344e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=8.4e-15 panw9=0 panw10=0 $X=121270 $Y=42830 $D=111
M8738 3910 3909 3912 VDD lppfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.77816e-13 as=1.52483e-13 pd=1.60444e-06 ps=1.35111e-06 nrd=0.307853 nrs=0.263993 sa=6.22105e-07 sb=9.05789e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=121750 $Y=42830 $D=111
M8739 3913 3912 3910 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9e-14 as=1.16984e-13 pd=8.6e-07 ps=1.05556e-06 nrd=0.36 nrs=0.467937 sa=5.896e-07 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=4.08e-14 panw10=0 $X=122230 $Y=43300 $D=111
M8740 3911 3914 3913 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.5e-13 as=9e-14 pd=1.1e-06 ps=8.6e-07 nrd=0.6 nrs=0.36 sa=1.0696e-06 sb=9.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=4.08e-14 panw10=0 $X=122710 $Y=43300 $D=111
M8741 VDD 403 3911 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.6e-13 as=1.5e-13 pd=1.71795e-06 ps=1.1e-06 nrd=0.64 nrs=0.6 sa=1.7608e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=4.08e-14 panw10=0 $X=123430 $Y=43300 $D=111
M8742 3915 3911 3912 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9e-14 as=1.6e-13 pd=8.6e-07 ps=1.64e-06 nrd=0.36 nrs=0.64 sa=3.2e-07 sb=7.856e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=124390 $Y=43040 $D=111
M8743 3914 403 3915 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.528e-13 as=9e-14 pd=1.64e-06 ps=8.6e-07 nrd=0.6112 nrs=0.36 sa=8e-07 sb=3.056e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=124870 $Y=43040 $D=111
M8744 VDD 3913 470 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=3.092e-13 pd=1.64e-06 ps=3.42e-06 nrd=0.140625 nrs=0.188721 sa=2.2625e-07 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=125690 $Y=42710 $D=111
M8745 845 3915 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=7.0625e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=126170 $Y=42710 $D=111
M8746 3917 189 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=40200 $Y=59650 $D=111
M8747 152 174 3917 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=40520 $Y=59650 $D=111
M8748 3918 174 152 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.512e-13 pd=1.08e-06 ps=1.2e-06 nrd=0.142857 nrs=0.214286 sa=1.12e-06 sb=1.96571e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=41000 $Y=59650 $D=111
M8749 VDD 189 3918 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.254e-13 as=1.008e-13 pd=1.57e-06 ps=1.08e-06 nrd=0.319444 nrs=0.142857 sa=1.48e-06 sb=1.94e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=41360 $Y=59650 $D=111
M8750 3919 180 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.254e-13 pd=1.04e-06 ps=1.57e-06 nrd=0.119048 nrs=0.319444 sa=2e-06 sb=1.41714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=41920 $Y=59650 $D=111
M8751 152 151 3919 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.572e-13 as=8.4e-14 pd=1.26e-06 ps=1.04e-06 nrd=0.222789 nrs=0.119048 sa=2e-06 sb=1.09714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=42240 $Y=59650 $D=111
M8752 3920 151 152 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.572e-13 pd=1.04e-06 ps=1.26e-06 nrd=0.119048 nrs=0.222789 sa=1.87714e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=42720 $Y=59590 $D=111
M8753 VDD 180 3920 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.675e-13 as=8.4e-14 pd=2.805e-06 ps=1.04e-06 nrd=0.520833 nrs=0.119048 sa=1.9e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=43040 $Y=59590 $D=111
M8754 3922 203 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=41400 $Y=21110 $D=111
M8755 173 182 3922 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=41720 $Y=21110 $D=111
M8756 3923 182 173 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.512e-13 pd=1.08e-06 ps=1.2e-06 nrd=0.142857 nrs=0.214286 sa=1.12e-06 sb=1.96571e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=42200 $Y=21110 $D=111
M8757 VDD 203 3923 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.254e-13 as=1.008e-13 pd=1.57e-06 ps=1.08e-06 nrd=0.319444 nrs=0.142857 sa=1.48e-06 sb=1.94e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=42560 $Y=21110 $D=111
M8758 3924 148 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.254e-13 pd=1.04e-06 ps=1.57e-06 nrd=0.119048 nrs=0.319444 sa=2e-06 sb=1.41714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=43120 $Y=21110 $D=111
M8759 173 165 3924 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.572e-13 as=8.4e-14 pd=1.26e-06 ps=1.04e-06 nrd=0.222789 nrs=0.119048 sa=2e-06 sb=1.09714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=43440 $Y=21110 $D=111
M8760 3925 165 173 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.572e-13 pd=1.04e-06 ps=1.26e-06 nrd=0.119048 nrs=0.222789 sa=1.87714e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=43920 $Y=21170 $D=111
M8761 VDD 148 3925 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.675e-13 as=8.4e-14 pd=2.805e-06 ps=1.04e-06 nrd=0.520833 nrs=0.119048 sa=1.9e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=44240 $Y=21170 $D=111
M8762 3927 179 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=43800 $Y=64310 $D=111
M8763 894 189 3927 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=44120 $Y=64310 $D=111
M8764 3928 189 894 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.512e-13 pd=1.08e-06 ps=1.2e-06 nrd=0.142857 nrs=0.214286 sa=1.12e-06 sb=1.96571e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=44600 $Y=64310 $D=111
M8765 VDD 179 3928 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.254e-13 as=1.008e-13 pd=1.57e-06 ps=1.08e-06 nrd=0.319444 nrs=0.142857 sa=1.48e-06 sb=1.94e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=44960 $Y=64310 $D=111
M8766 3929 174 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.254e-13 pd=1.04e-06 ps=1.57e-06 nrd=0.119048 nrs=0.319444 sa=2e-06 sb=1.41714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=45520 $Y=64310 $D=111
M8767 894 151 3929 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.572e-13 as=8.4e-14 pd=1.26e-06 ps=1.04e-06 nrd=0.222789 nrs=0.119048 sa=2e-06 sb=1.09714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=45840 $Y=64310 $D=111
M8768 3930 151 894 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.572e-13 pd=1.04e-06 ps=1.26e-06 nrd=0.119048 nrs=0.222789 sa=1.87714e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=46320 $Y=64370 $D=111
M8769 VDD 174 3930 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.675e-13 as=8.4e-14 pd=2.805e-06 ps=1.04e-06 nrd=0.520833 nrs=0.119048 sa=1.9e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=46640 $Y=64370 $D=111
M8770 3932 148 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=45400 $Y=42710 $D=111
M8771 812 185 3932 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=45720 $Y=42710 $D=111
M8772 3933 185 812 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.512e-13 pd=1.08e-06 ps=1.2e-06 nrd=0.142857 nrs=0.214286 sa=1.12e-06 sb=1.96571e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=46200 $Y=42710 $D=111
M8773 VDD 148 3933 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.254e-13 as=1.008e-13 pd=1.57e-06 ps=1.08e-06 nrd=0.319444 nrs=0.142857 sa=1.48e-06 sb=1.94e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=46560 $Y=42710 $D=111
M8774 3934 166 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.254e-13 pd=1.04e-06 ps=1.57e-06 nrd=0.119048 nrs=0.319444 sa=2e-06 sb=1.41714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=47120 $Y=42710 $D=111
M8775 812 168 3934 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.572e-13 as=8.4e-14 pd=1.26e-06 ps=1.04e-06 nrd=0.222789 nrs=0.119048 sa=2e-06 sb=1.09714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=47440 $Y=42710 $D=111
M8776 3935 168 812 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.572e-13 pd=1.04e-06 ps=1.26e-06 nrd=0.119048 nrs=0.222789 sa=1.87714e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=47920 $Y=42770 $D=111
M8777 VDD 166 3935 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.675e-13 as=8.4e-14 pd=2.805e-06 ps=1.04e-06 nrd=0.520833 nrs=0.119048 sa=1.9e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=48240 $Y=42770 $D=111
M8778 3937 148 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=51000 $Y=52450 $D=111
M8779 210 200 3937 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=51320 $Y=52450 $D=111
M8780 3938 200 210 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.512e-13 pd=1.08e-06 ps=1.2e-06 nrd=0.142857 nrs=0.214286 sa=1.12e-06 sb=1.96571e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=51800 $Y=52450 $D=111
M8781 VDD 148 3938 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.254e-13 as=1.008e-13 pd=1.57e-06 ps=1.08e-06 nrd=0.319444 nrs=0.142857 sa=1.48e-06 sb=1.94e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=52160 $Y=52450 $D=111
M8782 3939 185 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.254e-13 pd=1.04e-06 ps=1.57e-06 nrd=0.119048 nrs=0.319444 sa=2e-06 sb=1.41714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=52720 $Y=52450 $D=111
M8783 210 168 3939 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.572e-13 as=8.4e-14 pd=1.26e-06 ps=1.04e-06 nrd=0.222789 nrs=0.119048 sa=2e-06 sb=1.09714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=53040 $Y=52450 $D=111
M8784 3940 168 210 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.572e-13 pd=1.04e-06 ps=1.26e-06 nrd=0.119048 nrs=0.222789 sa=1.87714e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=53520 $Y=52390 $D=111
M8785 VDD 185 3940 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.675e-13 as=8.4e-14 pd=2.805e-06 ps=1.04e-06 nrd=0.520833 nrs=0.119048 sa=1.9e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=53840 $Y=52390 $D=111
M8786 3942 203 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=55000 $Y=28310 $D=111
M8787 227 148 3942 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=55320 $Y=28310 $D=111
M8788 3943 148 227 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.512e-13 pd=1.08e-06 ps=1.2e-06 nrd=0.142857 nrs=0.214286 sa=1.12e-06 sb=1.96571e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=55800 $Y=28310 $D=111
M8789 VDD 203 3943 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.254e-13 as=1.008e-13 pd=1.57e-06 ps=1.08e-06 nrd=0.319444 nrs=0.142857 sa=1.48e-06 sb=1.94e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=56160 $Y=28310 $D=111
M8790 3944 217 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.254e-13 pd=1.04e-06 ps=1.57e-06 nrd=0.119048 nrs=0.319444 sa=2e-06 sb=1.41714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=56720 $Y=28310 $D=111
M8791 227 198 3944 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.572e-13 as=8.4e-14 pd=1.26e-06 ps=1.04e-06 nrd=0.222789 nrs=0.119048 sa=2e-06 sb=1.09714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=57040 $Y=28310 $D=111
M8792 3945 198 227 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.572e-13 pd=1.04e-06 ps=1.26e-06 nrd=0.119048 nrs=0.222789 sa=1.87714e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=57520 $Y=28370 $D=111
M8793 VDD 217 3945 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.675e-13 as=8.4e-14 pd=2.805e-06 ps=1.04e-06 nrd=0.520833 nrs=0.119048 sa=1.9e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=57840 $Y=28370 $D=111
M8794 3947 291 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=67400 $Y=42710 $D=111
M8795 215 820 3947 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=67720 $Y=42710 $D=111
M8796 3948 820 215 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.512e-13 pd=1.08e-06 ps=1.2e-06 nrd=0.142857 nrs=0.214286 sa=1.12e-06 sb=1.96571e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=68200 $Y=42710 $D=111
M8797 VDD 291 3948 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.254e-13 as=1.008e-13 pd=1.57e-06 ps=1.08e-06 nrd=0.319444 nrs=0.142857 sa=1.48e-06 sb=1.94e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=68560 $Y=42710 $D=111
M8798 3949 267 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.254e-13 pd=1.04e-06 ps=1.57e-06 nrd=0.119048 nrs=0.319444 sa=2e-06 sb=1.41714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=69120 $Y=42710 $D=111
M8799 215 232 3949 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.572e-13 as=8.4e-14 pd=1.26e-06 ps=1.04e-06 nrd=0.222789 nrs=0.119048 sa=2e-06 sb=1.09714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=69440 $Y=42710 $D=111
M8800 3950 232 215 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.572e-13 pd=1.04e-06 ps=1.26e-06 nrd=0.119048 nrs=0.222789 sa=1.87714e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=69920 $Y=42770 $D=111
M8801 VDD 267 3950 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.675e-13 as=8.4e-14 pd=2.805e-06 ps=1.04e-06 nrd=0.520833 nrs=0.119048 sa=1.9e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=70240 $Y=42770 $D=111
M8802 3952 213 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=69000 $Y=57110 $D=111
M8803 266 280 3952 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=69320 $Y=57110 $D=111
M8804 3953 280 266 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.512e-13 pd=1.08e-06 ps=1.2e-06 nrd=0.142857 nrs=0.214286 sa=1.12e-06 sb=1.96571e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=69800 $Y=57110 $D=111
M8805 VDD 213 3953 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.254e-13 as=1.008e-13 pd=1.57e-06 ps=1.08e-06 nrd=0.319444 nrs=0.142857 sa=1.48e-06 sb=1.94e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=70160 $Y=57110 $D=111
M8806 3954 246 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.254e-13 pd=1.04e-06 ps=1.57e-06 nrd=0.119048 nrs=0.319444 sa=2e-06 sb=1.41714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=70720 $Y=57110 $D=111
M8807 266 255 3954 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.572e-13 as=8.4e-14 pd=1.26e-06 ps=1.04e-06 nrd=0.222789 nrs=0.119048 sa=2e-06 sb=1.09714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=71040 $Y=57110 $D=111
M8808 3955 255 266 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.572e-13 pd=1.04e-06 ps=1.26e-06 nrd=0.119048 nrs=0.222789 sa=1.87714e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=71520 $Y=57170 $D=111
M8809 VDD 246 3955 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.675e-13 as=8.4e-14 pd=2.805e-06 ps=1.04e-06 nrd=0.520833 nrs=0.119048 sa=1.9e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=71840 $Y=57170 $D=111
M8810 3957 319 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=87400 $Y=42710 $D=111
M8811 320 336 3957 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=87720 $Y=42710 $D=111
M8812 3958 336 320 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.512e-13 pd=1.08e-06 ps=1.2e-06 nrd=0.142857 nrs=0.214286 sa=1.12e-06 sb=1.96571e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=88200 $Y=42710 $D=111
M8813 VDD 319 3958 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.254e-13 as=1.008e-13 pd=1.57e-06 ps=1.08e-06 nrd=0.319444 nrs=0.142857 sa=1.48e-06 sb=1.94e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=88560 $Y=42710 $D=111
M8814 3959 313 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.254e-13 pd=1.04e-06 ps=1.57e-06 nrd=0.119048 nrs=0.319444 sa=2e-06 sb=1.41714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=89120 $Y=42710 $D=111
M8815 320 330 3959 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.572e-13 as=8.4e-14 pd=1.26e-06 ps=1.04e-06 nrd=0.222789 nrs=0.119048 sa=2e-06 sb=1.09714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=89440 $Y=42710 $D=111
M8816 3960 330 320 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.572e-13 pd=1.04e-06 ps=1.26e-06 nrd=0.119048 nrs=0.222789 sa=1.87714e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=89920 $Y=42770 $D=111
M8817 VDD 313 3960 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.675e-13 as=8.4e-14 pd=2.805e-06 ps=1.04e-06 nrd=0.520833 nrs=0.119048 sa=1.9e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=90240 $Y=42770 $D=111
M8818 3962 419 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.688e-13 pd=1.04e-06 ps=2.32e-06 nrd=0.119048 nrs=0.380952 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=114200 $Y=42710 $D=111
M8819 446 410 3962 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=114520 $Y=42710 $D=111
M8820 3963 410 446 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.512e-13 pd=1.08e-06 ps=1.2e-06 nrd=0.142857 nrs=0.214286 sa=1.12e-06 sb=1.96571e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=115000 $Y=42710 $D=111
M8821 VDD 419 3963 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.254e-13 as=1.008e-13 pd=1.57e-06 ps=1.08e-06 nrd=0.319444 nrs=0.142857 sa=1.48e-06 sb=1.94e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=115360 $Y=42710 $D=111
M8822 3964 400 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=2.254e-13 pd=1.04e-06 ps=1.57e-06 nrd=0.119048 nrs=0.319444 sa=2e-06 sb=1.41714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=115920 $Y=42710 $D=111
M8823 446 416 3964 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.572e-13 as=8.4e-14 pd=1.26e-06 ps=1.04e-06 nrd=0.222789 nrs=0.119048 sa=2e-06 sb=1.09714e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.68e-14 panw10=0 $X=116240 $Y=42710 $D=111
M8824 3965 416 446 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.572e-13 pd=1.04e-06 ps=1.26e-06 nrd=0.119048 nrs=0.222789 sa=1.87714e-06 sb=6.8e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=116720 $Y=42770 $D=111
M8825 VDD 400 3965 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.675e-13 as=8.4e-14 pd=2.805e-06 ps=1.04e-06 nrd=0.520833 nrs=0.119048 sa=1.9e-06 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=4.8e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.4e-14 panw10=0 $X=117040 $Y=42770 $D=111
M8826 3974 357 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=96060 $Y=45080 $D=111
M8827 3967 3969 3974 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=96380 $Y=45080 $D=111
M8828 VDD 329 3967 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.362e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73724 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=96860 $Y=45080 $D=111
M8829 VDD clk 3966 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.043e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15816 nrs=0.761905 sa=3.2e-07 sb=6.82857e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=97380 $Y=45670 $D=111
M8830 3969 3966 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.362e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73724 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=97890 $Y=45790 $D=111
M8831 3976 3966 3967 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=98450 $Y=45310 $D=111
M8832 VDD 3968 3976 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=98770 $Y=45310 $D=111
M8833 3968 3967 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=99310 $Y=45310 $D=111
M8834 3970 3966 3968 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=100140 $Y=45060 $D=111
M8835 3979 3969 3970 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=100870 $Y=45060 $D=111
M8836 VDD 3972 3979 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=101200 $Y=45060 $D=111
M8837 3972 329 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=101660 $Y=45130 $D=111
M8838 VDD 3970 3972 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.14961e-13 as=8.48e-14 pd=7.79363e-07 ps=1.01e-06 nrd=1.46633 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=102220 $Y=44840 $D=111
M8839 3971 3972 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.14961e-13 pd=1.2e-06 ps=7.79363e-07 nrd=1.14286 nrs=1.46633 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=102830 $Y=45480 $D=111
M8840 VDD 3971 942 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.62767e-13 as=2.048e-13 pd=1.7814e-06 ps=1.92e-06 nrd=0.641521 nrs=0.5 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=103770 $Y=45450 $D=111
M8841 359 3972 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.62767e-13 pd=1.92e-06 ps=1.7814e-06 nrd=0.5 nrs=0.641521 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=104270 $Y=45450 $D=111
M8842 3990 369 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=103260 $Y=57840 $D=111
M8843 3983 3985 3990 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=103580 $Y=57840 $D=111
M8844 VDD 374 3983 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.362e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73724 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=104060 $Y=57840 $D=111
M8845 VDD clk 3982 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.043e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15816 nrs=0.761905 sa=3.2e-07 sb=6.82857e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=104580 $Y=57110 $D=111
M8846 3985 3982 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.362e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73724 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=105090 $Y=57130 $D=111
M8847 3992 3982 3983 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=105650 $Y=57610 $D=111
M8848 VDD 3984 3992 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=105970 $Y=57610 $D=111
M8849 3984 3983 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=106510 $Y=57610 $D=111
M8850 3986 3982 3984 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=107340 $Y=57860 $D=111
M8851 3995 3985 3986 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=108070 $Y=57860 $D=111
M8852 VDD 3988 3995 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=108400 $Y=57860 $D=111
M8853 3988 374 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=108860 $Y=57790 $D=111
M8854 VDD 3986 3988 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.14961e-13 as=8.48e-14 pd=7.79363e-07 ps=1.01e-06 nrd=1.46633 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=109420 $Y=58080 $D=111
M8855 3987 3988 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.14961e-13 pd=1.2e-06 ps=7.79363e-07 nrd=1.14286 nrs=1.46633 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=110030 $Y=57440 $D=111
M8856 VDD 3987 837 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.62767e-13 as=2.048e-13 pd=1.7814e-06 ps=1.92e-06 nrd=0.641521 nrs=0.5 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=110970 $Y=57110 $D=111
M8857 418 3988 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.62767e-13 pd=1.92e-06 ps=1.7814e-06 nrd=0.5 nrs=0.641521 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=111470 $Y=57110 $D=111
M8858 4006 835 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=112060 $Y=52280 $D=111
M8859 3999 4001 4006 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=112380 $Y=52280 $D=111
M8860 VDD 425 3999 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.362e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73724 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=112860 $Y=52280 $D=111
M8861 VDD clk 3998 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.043e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15816 nrs=0.761905 sa=3.2e-07 sb=6.82857e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=113380 $Y=52870 $D=111
M8862 4001 3998 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.362e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73724 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=0 panw8=0 panw9=0 panw10=0 $X=113890 $Y=52990 $D=111
M8863 4008 3998 3999 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=114450 $Y=52510 $D=111
M8864 VDD 4000 4008 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=114770 $Y=52510 $D=111
M8865 4000 3999 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=115310 $Y=52510 $D=111
M8866 4002 3998 4000 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.65e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=116140 $Y=52260 $D=111
M8867 4011 4001 4002 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=9.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=116870 $Y=52260 $D=111
M8868 VDD 4004 4011 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.76667e-14 as=2.94e-14 pd=8.86667e-07 ps=4.9e-07 nrd=0.990646 nrs=0.375 sa=1.72321e-06 sb=5.9e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=117200 $Y=52260 $D=111
M8869 4004 425 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.48e-14 as=7.76667e-14 pd=1.01e-06 ps=8.86667e-07 nrd=1.08163 nrs=0.990646 sa=1.565e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-15 panw9=3.12e-14 panw10=0 $X=117660 $Y=52330 $D=111
M8870 VDD 4002 4004 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.14961e-13 as=8.48e-14 pd=7.79363e-07 ps=1.01e-06 nrd=1.46633 nrs=1.08163 sa=3.6e-07 sb=1.49e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.56e-14 panw10=1.8e-14 $X=118220 $Y=52040 $D=111
M8871 4003 4004 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.96e-14 as=1.14961e-13 pd=1.2e-06 ps=7.79363e-07 nrd=1.14286 nrs=1.46633 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=1.32e-14 panw9=0 panw10=0 $X=118830 $Y=52680 $D=111
M8872 VDD 4003 943 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.62767e-13 as=2.048e-13 pd=1.7814e-06 ps=1.92e-06 nrd=0.641521 nrs=0.5 sa=3.2e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=119770 $Y=52650 $D=111
M8873 452 4004 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.62767e-13 pd=1.92e-06 ps=1.7814e-06 nrd=0.5 nrs=0.641521 sa=8.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=120270 $Y=52650 $D=111
M8874 4015 93 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.1339e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=6.5e-14 panw8=8.14e-14 panw9=1.44e-14 panw10=0 $X=8810 $Y=23670 $D=111
M8875 VDD 93 4015 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9813e-13 as=1.476e-13 pd=1.89486e-06 ps=1.18e-06 nrd=0.294661 nrs=0.219512 sa=8e-07 sb=6.53902e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.128e-13 panw10=0 $X=9290 $Y=23670 $D=111
M8876 4014 93 VDD VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.074e-13 as=1.5947e-13 pd=1.96e-06 ps=1.52514e-06 nrd=0.476125 nrs=0.366093 sa=1.24e-06 sb=3.14242e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=7.92e-14 $X=9730 $Y=23830 $D=111
M8877 VDD 4014 4016 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.104e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.312909 sa=2.56585e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=10570 $Y=23340 $D=111
M8878 4016 4014 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=7.36585e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=11050 $Y=23340 $D=111
M8879 4017 4018 4016 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.21659e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=11530 $Y=23340 $D=111
M8880 4016 4018 4017 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.69659e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=12010 $Y=23340 $D=111
M8881 4017 90 4015 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.69463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=12950 $Y=23660 $D=111
M8882 4015 90 4017 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=8e-07 sb=1.21463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=13430 $Y=23660 $D=111
M8883 4020 4018 4015 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.28e-06 sb=7.34634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=13910 $Y=23660 $D=111
M8884 4015 4018 4020 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.088e-13 as=1.476e-13 pd=2.36e-06 ps=1.18e-06 nrd=0.310529 nrs=0.219512 sa=1.76e-06 sb=2.54634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=14390 $Y=23660 $D=111
M8885 4020 90 4016 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=3.176e-13 pd=1.18e-06 ps=2.68e-06 nrd=0.219512 nrs=0.472338 sa=3.32683e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=15250 $Y=23340 $D=111
M8886 4016 90 4020 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.4e-13 as=1.476e-13 pd=2.68e-06 ps=1.18e-06 nrd=0.505651 nrs=0.219512 sa=8.12683e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=15730 $Y=23340 $D=111
M8887 VDD 90 4018 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.339e-13 as=3.392e-13 pd=1.69e-06 ps=2.76e-06 nrd=0.29717 nrs=0.301887 sa=3.2e-07 sb=1.91406e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=16790 $Y=23190 $D=111
M8888 4018 90 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.74673e-13 as=3.339e-13 pd=1.84713e-06 ps=1.69e-06 nrd=0.333458 nrs=0.29717 sa=1.07e-06 sb=1.60358e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=17540 $Y=23190 $D=111
M8889 4019 4020 4018 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93608e-13 as=3.39327e-13 pd=1.82905e-06 ps=1.67287e-06 nrd=0.318586 nrs=0.368193 sa=1.86635e-06 sb=1.42469e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=18350 $Y=23180 $D=111
M8890 4022 4017 4019 VDD lppfet w=9.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.20041e-13 as=2.87492e-13 pd=1.66774e-06 ps=1.79095e-06 nrd=0.249028 nrs=0.325364 sa=1.44926e-06 sb=1.38872e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=19010 $Y=23510 $D=111
M8891 4023 4020 4022 VDD lppfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.78404e-13 as=2.15359e-13 pd=1.40371e-06 ps=1.63226e-06 nrd=0.21078 nrs=0.254441 sa=1.4087e-06 sb=1.70522e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=19520 $Y=23190 $D=111
M8892 4021 4017 4023 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.244e-13 as=1.97796e-13 pd=1.46e-06 ps=1.55629e-06 nrd=0.215686 nrs=0.190115 sa=1.39961e-06 sb=1.41e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=20000 $Y=23290 $D=111
M8893 VDD 4022 4021 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.33972e-13 as=2.244e-13 pd=1.57708e-06 ps=1.46e-06 nrd=0.224887 nrs=0.215686 sa=1.6302e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=20560 $Y=23290 $D=111
M8894 4022 66 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.764e-13 as=2.982e-13 pd=3.24e-06 ps=2.01e-06 nrd=0.222722 nrs=0.17645 sa=1.51538e-06 sb=2.89538e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=21120 $Y=23190 $D=111
M8895 VDD 4019 17 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.054e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.247437 sa=3.16719e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=22160 $Y=23210 $D=111
M8896 39 4023 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.352e-13 as=2.304e-13 pd=3.24e-06 ps=1.64e-06 nrd=0.265625 nrs=0.140625 sa=7.96719e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=22640 $Y=23210 $D=111
M8897 4025 150 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.1339e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=6.5e-14 panw8=8.14e-14 panw9=1.44e-14 panw10=0 $X=8810 $Y=42710 $D=111
M8898 VDD 150 4025 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9813e-13 as=1.476e-13 pd=1.89486e-06 ps=1.18e-06 nrd=0.294661 nrs=0.219512 sa=8e-07 sb=6.53902e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.128e-13 panw10=0 $X=9290 $Y=42710 $D=111
M8899 4024 150 VDD VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.074e-13 as=1.5947e-13 pd=1.96e-06 ps=1.52514e-06 nrd=0.476125 nrs=0.366093 sa=1.24e-06 sb=3.14242e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=7.92e-14 $X=9730 $Y=42710 $D=111
M8900 VDD 4024 4026 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.104e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.312909 sa=2.56585e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=10570 $Y=43040 $D=111
M8901 4026 4024 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=7.36585e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=11050 $Y=43040 $D=111
M8902 4027 4028 4026 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.21659e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=11530 $Y=43040 $D=111
M8903 4026 4028 4027 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.69659e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=12010 $Y=43040 $D=111
M8904 4027 53 4025 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.69463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=12950 $Y=42720 $D=111
M8905 4025 53 4027 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=8e-07 sb=1.21463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=13430 $Y=42720 $D=111
M8906 4030 4028 4025 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.28e-06 sb=7.34634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=13910 $Y=42720 $D=111
M8907 4025 4028 4030 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.088e-13 as=1.476e-13 pd=2.36e-06 ps=1.18e-06 nrd=0.310529 nrs=0.219512 sa=1.76e-06 sb=2.54634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=14390 $Y=42720 $D=111
M8908 4030 53 4026 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=3.176e-13 pd=1.18e-06 ps=2.68e-06 nrd=0.219512 nrs=0.472338 sa=3.32683e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=15250 $Y=43040 $D=111
M8909 4026 53 4030 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.4e-13 as=1.476e-13 pd=2.68e-06 ps=1.18e-06 nrd=0.505651 nrs=0.219512 sa=8.12683e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=15730 $Y=43040 $D=111
M8910 VDD 53 4028 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.339e-13 as=3.392e-13 pd=1.69e-06 ps=2.76e-06 nrd=0.29717 nrs=0.301887 sa=3.2e-07 sb=1.91406e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=16790 $Y=42950 $D=111
M8911 4028 53 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.74673e-13 as=3.339e-13 pd=1.84713e-06 ps=1.69e-06 nrd=0.333458 nrs=0.29717 sa=1.07e-06 sb=1.60358e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=17540 $Y=42950 $D=111
M8912 4029 4030 4028 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93608e-13 as=3.39327e-13 pd=1.82905e-06 ps=1.67287e-06 nrd=0.318586 nrs=0.368193 sa=1.86635e-06 sb=1.42469e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=18350 $Y=43060 $D=111
M8913 4032 4027 4029 VDD lppfet w=9.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.20041e-13 as=2.87492e-13 pd=1.66774e-06 ps=1.79095e-06 nrd=0.249028 nrs=0.325364 sa=1.44926e-06 sb=1.38872e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=19010 $Y=42750 $D=111
M8914 4033 4030 4032 VDD lppfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.78404e-13 as=2.15359e-13 pd=1.40371e-06 ps=1.63226e-06 nrd=0.21078 nrs=0.254441 sa=1.4087e-06 sb=1.70522e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=19520 $Y=43090 $D=111
M8915 4031 4027 4033 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.244e-13 as=1.97796e-13 pd=1.46e-06 ps=1.55629e-06 nrd=0.215686 nrs=0.190115 sa=1.39961e-06 sb=1.41e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=20000 $Y=42890 $D=111
M8916 VDD 4032 4031 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.33972e-13 as=2.244e-13 pd=1.57708e-06 ps=1.46e-06 nrd=0.224887 nrs=0.215686 sa=1.6302e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=20560 $Y=42890 $D=111
M8917 4032 94 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.764e-13 as=2.982e-13 pd=3.24e-06 ps=2.01e-06 nrd=0.222722 nrs=0.17645 sa=1.51538e-06 sb=2.89538e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=21120 $Y=42710 $D=111
M8918 VDD 4029 944 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.054e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.247437 sa=3.16719e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=22160 $Y=42710 $D=111
M8919 8 4033 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.352e-13 as=2.304e-13 pd=3.24e-06 ps=1.64e-06 nrd=0.265625 nrs=0.140625 sa=7.96719e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=22640 $Y=42710 $D=111
M8920 4035 92 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.1339e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=22010 $Y=49910 $D=111
M8921 VDD 92 4035 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9813e-13 as=1.476e-13 pd=1.89486e-06 ps=1.18e-06 nrd=0.294661 nrs=0.219512 sa=8e-07 sb=6.53902e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=22490 $Y=49910 $D=111
M8922 4034 92 VDD VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.074e-13 as=1.5947e-13 pd=1.96e-06 ps=1.52514e-06 nrd=0.476125 nrs=0.366093 sa=1.24e-06 sb=3.14242e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=22930 $Y=49910 $D=111
M8923 VDD 4034 4036 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.104e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.312909 sa=2.56585e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=23770 $Y=50240 $D=111
M8924 4036 4034 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=7.36585e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=24250 $Y=50240 $D=111
M8925 4037 4038 4036 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.21659e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=24730 $Y=50240 $D=111
M8926 4036 4038 4037 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.69659e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=25210 $Y=50240 $D=111
M8927 4037 120 4035 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.69463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=26150 $Y=49920 $D=111
M8928 4035 120 4037 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=8e-07 sb=1.21463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=26630 $Y=49920 $D=111
M8929 4040 4038 4035 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.28e-06 sb=7.34634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=27110 $Y=49920 $D=111
M8930 4035 4038 4040 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.088e-13 as=1.476e-13 pd=2.36e-06 ps=1.18e-06 nrd=0.310529 nrs=0.219512 sa=1.76e-06 sb=2.54634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=27590 $Y=49920 $D=111
M8931 4040 120 4036 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=3.176e-13 pd=1.18e-06 ps=2.68e-06 nrd=0.219512 nrs=0.472338 sa=3.32683e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=28450 $Y=50240 $D=111
M8932 4036 120 4040 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.4e-13 as=1.476e-13 pd=2.68e-06 ps=1.18e-06 nrd=0.505651 nrs=0.219512 sa=8.12683e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=28930 $Y=50240 $D=111
M8933 VDD 120 4038 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.339e-13 as=3.392e-13 pd=1.69e-06 ps=2.76e-06 nrd=0.29717 nrs=0.301887 sa=3.2e-07 sb=1.91406e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=29990 $Y=50150 $D=111
M8934 4038 120 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.74673e-13 as=3.339e-13 pd=1.84713e-06 ps=1.69e-06 nrd=0.333458 nrs=0.29717 sa=1.07e-06 sb=1.60358e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=30740 $Y=50150 $D=111
M8935 4039 4040 4038 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93608e-13 as=3.39327e-13 pd=1.82905e-06 ps=1.67287e-06 nrd=0.318586 nrs=0.368193 sa=1.86635e-06 sb=1.42469e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=31550 $Y=50260 $D=111
M8936 4042 4037 4039 VDD lppfet w=9.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.20041e-13 as=2.87492e-13 pd=1.66774e-06 ps=1.79095e-06 nrd=0.249028 nrs=0.325364 sa=1.44926e-06 sb=1.38872e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=32210 $Y=49950 $D=111
M8937 4043 4040 4042 VDD lppfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.78404e-13 as=2.15359e-13 pd=1.40371e-06 ps=1.63226e-06 nrd=0.21078 nrs=0.254441 sa=1.4087e-06 sb=1.70522e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=32720 $Y=50290 $D=111
M8938 4041 4037 4043 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.244e-13 as=1.97796e-13 pd=1.46e-06 ps=1.55629e-06 nrd=0.215686 nrs=0.190115 sa=1.39961e-06 sb=1.41e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=33200 $Y=50090 $D=111
M8939 VDD 4042 4041 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.33972e-13 as=2.244e-13 pd=1.57708e-06 ps=1.46e-06 nrd=0.224887 nrs=0.215686 sa=1.6302e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=33760 $Y=50090 $D=111
M8940 4042 197 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.764e-13 as=2.982e-13 pd=3.24e-06 ps=2.01e-06 nrd=0.222722 nrs=0.17645 sa=1.51538e-06 sb=2.89538e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=34320 $Y=49910 $D=111
M8941 VDD 4039 121 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.054e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.247437 sa=3.16719e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=35360 $Y=49910 $D=111
M8942 124 4043 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.352e-13 as=2.304e-13 pd=3.24e-06 ps=1.64e-06 nrd=0.265625 nrs=0.140625 sa=7.96719e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=35840 $Y=49910 $D=111
M8943 4045 77 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.1339e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=23610 $Y=23670 $D=111
M8944 VDD 77 4045 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9813e-13 as=1.476e-13 pd=1.89486e-06 ps=1.18e-06 nrd=0.294661 nrs=0.219512 sa=8e-07 sb=6.53902e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=24090 $Y=23670 $D=111
M8945 4044 77 VDD VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.074e-13 as=1.5947e-13 pd=1.96e-06 ps=1.52514e-06 nrd=0.476125 nrs=0.366093 sa=1.24e-06 sb=3.14242e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=24530 $Y=23830 $D=111
M8946 VDD 4044 4046 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.104e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.312909 sa=2.56585e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=25370 $Y=23340 $D=111
M8947 4046 4044 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=7.36585e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=25850 $Y=23340 $D=111
M8948 4047 4048 4046 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.21659e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=26330 $Y=23340 $D=111
M8949 4046 4048 4047 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.69659e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=26810 $Y=23340 $D=111
M8950 4047 155 4045 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.69463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=27750 $Y=23660 $D=111
M8951 4045 155 4047 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=8e-07 sb=1.21463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=28230 $Y=23660 $D=111
M8952 4050 4048 4045 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.28e-06 sb=7.34634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=28710 $Y=23660 $D=111
M8953 4045 4048 4050 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.088e-13 as=1.476e-13 pd=2.36e-06 ps=1.18e-06 nrd=0.310529 nrs=0.219512 sa=1.76e-06 sb=2.54634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=29190 $Y=23660 $D=111
M8954 4050 155 4046 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=3.176e-13 pd=1.18e-06 ps=2.68e-06 nrd=0.219512 nrs=0.472338 sa=3.32683e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=30050 $Y=23340 $D=111
M8955 4046 155 4050 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.4e-13 as=1.476e-13 pd=2.68e-06 ps=1.18e-06 nrd=0.505651 nrs=0.219512 sa=8.12683e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=30530 $Y=23340 $D=111
M8956 VDD 155 4048 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.339e-13 as=3.392e-13 pd=1.69e-06 ps=2.76e-06 nrd=0.29717 nrs=0.301887 sa=3.2e-07 sb=1.91406e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=31590 $Y=23190 $D=111
M8957 4048 155 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.74673e-13 as=3.339e-13 pd=1.84713e-06 ps=1.69e-06 nrd=0.333458 nrs=0.29717 sa=1.07e-06 sb=1.60358e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=32340 $Y=23190 $D=111
M8958 4049 4050 4048 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93608e-13 as=3.39327e-13 pd=1.82905e-06 ps=1.67287e-06 nrd=0.318586 nrs=0.368193 sa=1.86635e-06 sb=1.42469e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=33150 $Y=23180 $D=111
M8959 4052 4047 4049 VDD lppfet w=9.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.20041e-13 as=2.87492e-13 pd=1.66774e-06 ps=1.79095e-06 nrd=0.249028 nrs=0.325364 sa=1.44926e-06 sb=1.38872e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=33810 $Y=23510 $D=111
M8960 4053 4050 4052 VDD lppfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.78404e-13 as=2.15359e-13 pd=1.40371e-06 ps=1.63226e-06 nrd=0.21078 nrs=0.254441 sa=1.4087e-06 sb=1.70522e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=34320 $Y=23190 $D=111
M8961 4051 4047 4053 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.244e-13 as=1.97796e-13 pd=1.46e-06 ps=1.55629e-06 nrd=0.215686 nrs=0.190115 sa=1.39961e-06 sb=1.41e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=34800 $Y=23290 $D=111
M8962 VDD 4052 4051 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.33972e-13 as=2.244e-13 pd=1.57708e-06 ps=1.46e-06 nrd=0.224887 nrs=0.215686 sa=1.6302e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=35360 $Y=23290 $D=111
M8963 4052 126 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.764e-13 as=2.982e-13 pd=3.24e-06 ps=2.01e-06 nrd=0.222722 nrs=0.17645 sa=1.51538e-06 sb=2.89538e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=35920 $Y=23190 $D=111
M8964 VDD 4049 133 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.054e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.247437 sa=3.16719e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=36960 $Y=23210 $D=111
M8965 130 4053 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.352e-13 as=2.304e-13 pd=3.24e-06 ps=1.64e-06 nrd=0.265625 nrs=0.140625 sa=7.96719e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=37440 $Y=23210 $D=111
M8966 4055 149 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.1339e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=38810 $Y=71510 $D=111
M8967 VDD 149 4055 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9813e-13 as=1.476e-13 pd=1.89486e-06 ps=1.18e-06 nrd=0.294661 nrs=0.219512 sa=8e-07 sb=6.53902e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=39290 $Y=71510 $D=111
M8968 4054 149 VDD VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.074e-13 as=1.5947e-13 pd=1.96e-06 ps=1.52514e-06 nrd=0.476125 nrs=0.366093 sa=1.24e-06 sb=3.14242e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=39730 $Y=71510 $D=111
M8969 VDD 4054 4056 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.104e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.312909 sa=2.56585e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=40570 $Y=71840 $D=111
M8970 4056 4054 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=7.36585e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=41050 $Y=71840 $D=111
M8971 4057 4058 4056 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.21659e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=41530 $Y=71840 $D=111
M8972 4056 4058 4057 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.69659e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=42010 $Y=71840 $D=111
M8973 4057 225 4055 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.69463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=42950 $Y=71520 $D=111
M8974 4055 225 4057 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=8e-07 sb=1.21463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=43430 $Y=71520 $D=111
M8975 4060 4058 4055 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.28e-06 sb=7.34634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=43910 $Y=71520 $D=111
M8976 4055 4058 4060 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.088e-13 as=1.476e-13 pd=2.36e-06 ps=1.18e-06 nrd=0.310529 nrs=0.219512 sa=1.76e-06 sb=2.54634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=44390 $Y=71520 $D=111
M8977 4060 225 4056 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=3.176e-13 pd=1.18e-06 ps=2.68e-06 nrd=0.219512 nrs=0.472338 sa=3.32683e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=45250 $Y=71840 $D=111
M8978 4056 225 4060 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.4e-13 as=1.476e-13 pd=2.68e-06 ps=1.18e-06 nrd=0.505651 nrs=0.219512 sa=8.12683e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=45730 $Y=71840 $D=111
M8979 VDD 225 4058 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.339e-13 as=3.392e-13 pd=1.69e-06 ps=2.76e-06 nrd=0.29717 nrs=0.301887 sa=3.2e-07 sb=1.91406e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=46790 $Y=71750 $D=111
M8980 4058 225 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.74673e-13 as=3.339e-13 pd=1.84713e-06 ps=1.69e-06 nrd=0.333458 nrs=0.29717 sa=1.07e-06 sb=1.60358e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=47540 $Y=71750 $D=111
M8981 4059 4060 4058 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93608e-13 as=3.39327e-13 pd=1.82905e-06 ps=1.67287e-06 nrd=0.318586 nrs=0.368193 sa=1.86635e-06 sb=1.42469e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=48350 $Y=71860 $D=111
M8982 4062 4057 4059 VDD lppfet w=9.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.20041e-13 as=2.87492e-13 pd=1.66774e-06 ps=1.79095e-06 nrd=0.249028 nrs=0.325364 sa=1.44926e-06 sb=1.38872e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=49010 $Y=71550 $D=111
M8983 4063 4060 4062 VDD lppfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.78404e-13 as=2.15359e-13 pd=1.40371e-06 ps=1.63226e-06 nrd=0.21078 nrs=0.254441 sa=1.4087e-06 sb=1.70522e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=49520 $Y=71890 $D=111
M8984 4061 4057 4063 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.244e-13 as=1.97796e-13 pd=1.46e-06 ps=1.55629e-06 nrd=0.215686 nrs=0.190115 sa=1.39961e-06 sb=1.41e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=50000 $Y=71690 $D=111
M8985 VDD 4062 4061 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.33972e-13 as=2.244e-13 pd=1.57708e-06 ps=1.46e-06 nrd=0.224887 nrs=0.215686 sa=1.6302e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=50560 $Y=71690 $D=111
M8986 4062 196 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.764e-13 as=2.982e-13 pd=3.24e-06 ps=2.01e-06 nrd=0.222722 nrs=0.17645 sa=1.51538e-06 sb=2.89538e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=51120 $Y=71510 $D=111
M8987 VDD 4059 191 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.054e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.247437 sa=3.16719e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=52160 $Y=71510 $D=111
M8988 69 4063 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.352e-13 as=2.304e-13 pd=3.24e-06 ps=1.64e-06 nrd=0.265625 nrs=0.140625 sa=7.96719e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=52640 $Y=71510 $D=111
M8989 4065 152 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.1339e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=39210 $Y=66870 $D=111
M8990 VDD 152 4065 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9813e-13 as=1.476e-13 pd=1.89486e-06 ps=1.18e-06 nrd=0.294661 nrs=0.219512 sa=8e-07 sb=6.53902e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=39690 $Y=66870 $D=111
M8991 4064 152 VDD VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.074e-13 as=1.5947e-13 pd=1.96e-06 ps=1.52514e-06 nrd=0.476125 nrs=0.366093 sa=1.24e-06 sb=3.14242e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=40130 $Y=67030 $D=111
M8992 VDD 4064 4066 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.104e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.312909 sa=2.56585e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=40970 $Y=66540 $D=111
M8993 4066 4064 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=7.36585e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=41450 $Y=66540 $D=111
M8994 4067 4068 4066 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.21659e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=41930 $Y=66540 $D=111
M8995 4066 4068 4067 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.69659e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=42410 $Y=66540 $D=111
M8996 4067 250 4065 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.69463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=43350 $Y=66860 $D=111
M8997 4065 250 4067 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=8e-07 sb=1.21463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=43830 $Y=66860 $D=111
M8998 4070 4068 4065 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.28e-06 sb=7.34634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=44310 $Y=66860 $D=111
M8999 4065 4068 4070 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.088e-13 as=1.476e-13 pd=2.36e-06 ps=1.18e-06 nrd=0.310529 nrs=0.219512 sa=1.76e-06 sb=2.54634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=44790 $Y=66860 $D=111
M9000 4070 250 4066 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=3.176e-13 pd=1.18e-06 ps=2.68e-06 nrd=0.219512 nrs=0.472338 sa=3.32683e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=45650 $Y=66540 $D=111
M9001 4066 250 4070 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.4e-13 as=1.476e-13 pd=2.68e-06 ps=1.18e-06 nrd=0.505651 nrs=0.219512 sa=8.12683e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=46130 $Y=66540 $D=111
M9002 VDD 250 4068 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.339e-13 as=3.392e-13 pd=1.69e-06 ps=2.76e-06 nrd=0.29717 nrs=0.301887 sa=3.2e-07 sb=1.91406e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=47190 $Y=66390 $D=111
M9003 4068 250 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.74673e-13 as=3.339e-13 pd=1.84713e-06 ps=1.69e-06 nrd=0.333458 nrs=0.29717 sa=1.07e-06 sb=1.60358e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=47940 $Y=66390 $D=111
M9004 4069 4070 4068 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93608e-13 as=3.39327e-13 pd=1.82905e-06 ps=1.67287e-06 nrd=0.318586 nrs=0.368193 sa=1.86635e-06 sb=1.42469e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=48750 $Y=66380 $D=111
M9005 4072 4067 4069 VDD lppfet w=9.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.20041e-13 as=2.87492e-13 pd=1.66774e-06 ps=1.79095e-06 nrd=0.249028 nrs=0.325364 sa=1.44926e-06 sb=1.38872e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=49410 $Y=66710 $D=111
M9006 4073 4070 4072 VDD lppfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.78404e-13 as=2.15359e-13 pd=1.40371e-06 ps=1.63226e-06 nrd=0.21078 nrs=0.254441 sa=1.4087e-06 sb=1.70522e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=49920 $Y=66390 $D=111
M9007 4071 4067 4073 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.244e-13 as=1.97796e-13 pd=1.46e-06 ps=1.55629e-06 nrd=0.215686 nrs=0.190115 sa=1.39961e-06 sb=1.41e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=50400 $Y=66490 $D=111
M9008 VDD 4072 4071 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.33972e-13 as=2.244e-13 pd=1.57708e-06 ps=1.46e-06 nrd=0.224887 nrs=0.215686 sa=1.6302e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=50960 $Y=66490 $D=111
M9009 4072 190 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.764e-13 as=2.982e-13 pd=3.24e-06 ps=2.01e-06 nrd=0.222722 nrs=0.17645 sa=1.51538e-06 sb=2.89538e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=51520 $Y=66390 $D=111
M9010 VDD 4069 268 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.054e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.247437 sa=3.16719e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=52560 $Y=66410 $D=111
M9011 196 4073 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.352e-13 as=2.304e-13 pd=3.24e-06 ps=1.64e-06 nrd=0.265625 nrs=0.140625 sa=7.96719e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=53040 $Y=66410 $D=111
M9012 4075 279 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.1339e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=40810 $Y=45270 $D=111
M9013 VDD 279 4075 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9813e-13 as=1.476e-13 pd=1.89486e-06 ps=1.18e-06 nrd=0.294661 nrs=0.219512 sa=8e-07 sb=6.53902e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=41290 $Y=45270 $D=111
M9014 4074 279 VDD VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.074e-13 as=1.5947e-13 pd=1.96e-06 ps=1.52514e-06 nrd=0.476125 nrs=0.366093 sa=1.24e-06 sb=3.14242e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=41730 $Y=45430 $D=111
M9015 VDD 4074 4076 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.104e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.312909 sa=2.56585e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=42570 $Y=44940 $D=111
M9016 4076 4074 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=7.36585e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=43050 $Y=44940 $D=111
M9017 4077 4078 4076 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.21659e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=43530 $Y=44940 $D=111
M9018 4076 4078 4077 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.69659e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=44010 $Y=44940 $D=111
M9019 4077 812 4075 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.69463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=44950 $Y=45260 $D=111
M9020 4075 812 4077 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=8e-07 sb=1.21463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=45430 $Y=45260 $D=111
M9021 4080 4078 4075 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.28e-06 sb=7.34634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=45910 $Y=45260 $D=111
M9022 4075 4078 4080 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.088e-13 as=1.476e-13 pd=2.36e-06 ps=1.18e-06 nrd=0.310529 nrs=0.219512 sa=1.76e-06 sb=2.54634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=46390 $Y=45260 $D=111
M9023 4080 812 4076 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=3.176e-13 pd=1.18e-06 ps=2.68e-06 nrd=0.219512 nrs=0.472338 sa=3.32683e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=47250 $Y=44940 $D=111
M9024 4076 812 4080 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.4e-13 as=1.476e-13 pd=2.68e-06 ps=1.18e-06 nrd=0.505651 nrs=0.219512 sa=8.12683e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=47730 $Y=44940 $D=111
M9025 VDD 812 4078 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.339e-13 as=3.392e-13 pd=1.69e-06 ps=2.76e-06 nrd=0.29717 nrs=0.301887 sa=3.2e-07 sb=1.91406e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=48790 $Y=44790 $D=111
M9026 4078 812 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.74673e-13 as=3.339e-13 pd=1.84713e-06 ps=1.69e-06 nrd=0.333458 nrs=0.29717 sa=1.07e-06 sb=1.60358e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=49540 $Y=44790 $D=111
M9027 4079 4080 4078 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93608e-13 as=3.39327e-13 pd=1.82905e-06 ps=1.67287e-06 nrd=0.318586 nrs=0.368193 sa=1.86635e-06 sb=1.42469e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=50350 $Y=44780 $D=111
M9028 4082 4077 4079 VDD lppfet w=9.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.20041e-13 as=2.87492e-13 pd=1.66774e-06 ps=1.79095e-06 nrd=0.249028 nrs=0.325364 sa=1.44926e-06 sb=1.38872e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=51010 $Y=45110 $D=111
M9029 4083 4080 4082 VDD lppfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.78404e-13 as=2.15359e-13 pd=1.40371e-06 ps=1.63226e-06 nrd=0.21078 nrs=0.254441 sa=1.4087e-06 sb=1.70522e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=51520 $Y=44790 $D=111
M9030 4081 4077 4083 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.244e-13 as=1.97796e-13 pd=1.46e-06 ps=1.55629e-06 nrd=0.215686 nrs=0.190115 sa=1.39961e-06 sb=1.41e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=52000 $Y=44890 $D=111
M9031 VDD 4082 4081 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.33972e-13 as=2.244e-13 pd=1.57708e-06 ps=1.46e-06 nrd=0.224887 nrs=0.215686 sa=1.6302e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=52560 $Y=44890 $D=111
M9032 4082 223 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.764e-13 as=2.982e-13 pd=3.24e-06 ps=2.01e-06 nrd=0.222722 nrs=0.17645 sa=1.51538e-06 sb=2.89538e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=53120 $Y=44790 $D=111
M9033 VDD 4079 149 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.054e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.247437 sa=3.16719e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=54160 $Y=44810 $D=111
M9034 197 4083 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.352e-13 as=2.304e-13 pd=3.24e-06 ps=1.64e-06 nrd=0.265625 nrs=0.140625 sa=7.96719e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=54640 $Y=44810 $D=111
M9035 4085 331 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.1339e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=84010 $Y=49910 $D=111
M9036 VDD 331 4085 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9813e-13 as=1.476e-13 pd=1.89486e-06 ps=1.18e-06 nrd=0.294661 nrs=0.219512 sa=8e-07 sb=6.53902e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=84490 $Y=49910 $D=111
M9037 4084 331 VDD VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.074e-13 as=1.5947e-13 pd=1.96e-06 ps=1.52514e-06 nrd=0.476125 nrs=0.366093 sa=1.24e-06 sb=3.14242e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=84930 $Y=49910 $D=111
M9038 VDD 4084 4086 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.104e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.312909 sa=2.56585e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=85770 $Y=50240 $D=111
M9039 4086 4084 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=7.36585e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=86250 $Y=50240 $D=111
M9040 4087 4088 4086 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.21659e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=86730 $Y=50240 $D=111
M9041 4086 4088 4087 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.69659e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=87210 $Y=50240 $D=111
M9042 4087 340 4085 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.69463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=88150 $Y=49920 $D=111
M9043 4085 340 4087 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=8e-07 sb=1.21463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=88630 $Y=49920 $D=111
M9044 4090 4088 4085 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.28e-06 sb=7.34634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=89110 $Y=49920 $D=111
M9045 4085 4088 4090 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.088e-13 as=1.476e-13 pd=2.36e-06 ps=1.18e-06 nrd=0.310529 nrs=0.219512 sa=1.76e-06 sb=2.54634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=89590 $Y=49920 $D=111
M9046 4090 340 4086 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=3.176e-13 pd=1.18e-06 ps=2.68e-06 nrd=0.219512 nrs=0.472338 sa=3.32683e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=90450 $Y=50240 $D=111
M9047 4086 340 4090 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.4e-13 as=1.476e-13 pd=2.68e-06 ps=1.18e-06 nrd=0.505651 nrs=0.219512 sa=8.12683e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=90930 $Y=50240 $D=111
M9048 VDD 340 4088 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.339e-13 as=3.392e-13 pd=1.69e-06 ps=2.76e-06 nrd=0.29717 nrs=0.301887 sa=3.2e-07 sb=1.91406e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=91990 $Y=50150 $D=111
M9049 4088 340 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.74673e-13 as=3.339e-13 pd=1.84713e-06 ps=1.69e-06 nrd=0.333458 nrs=0.29717 sa=1.07e-06 sb=1.60358e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=92740 $Y=50150 $D=111
M9050 4089 4090 4088 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93608e-13 as=3.39327e-13 pd=1.82905e-06 ps=1.67287e-06 nrd=0.318586 nrs=0.368193 sa=1.86635e-06 sb=1.42469e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=93550 $Y=50260 $D=111
M9051 4092 4087 4089 VDD lppfet w=9.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.20041e-13 as=2.87492e-13 pd=1.66774e-06 ps=1.79095e-06 nrd=0.249028 nrs=0.325364 sa=1.44926e-06 sb=1.38872e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=94210 $Y=49950 $D=111
M9052 4093 4090 4092 VDD lppfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.78404e-13 as=2.15359e-13 pd=1.40371e-06 ps=1.63226e-06 nrd=0.21078 nrs=0.254441 sa=1.4087e-06 sb=1.70522e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=94720 $Y=50290 $D=111
M9053 4091 4087 4093 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.244e-13 as=1.97796e-13 pd=1.46e-06 ps=1.55629e-06 nrd=0.215686 nrs=0.190115 sa=1.39961e-06 sb=1.41e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=95200 $Y=50090 $D=111
M9054 VDD 4092 4091 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.33972e-13 as=2.244e-13 pd=1.57708e-06 ps=1.46e-06 nrd=0.224887 nrs=0.215686 sa=1.6302e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=95760 $Y=50090 $D=111
M9055 4092 355 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.764e-13 as=2.982e-13 pd=3.24e-06 ps=2.01e-06 nrd=0.222722 nrs=0.17645 sa=1.51538e-06 sb=2.89538e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=96320 $Y=49910 $D=111
M9056 VDD 4089 381 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.054e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.247437 sa=3.16719e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=97360 $Y=49910 $D=111
M9057 831 4093 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.352e-13 as=2.304e-13 pd=3.24e-06 ps=1.64e-06 nrd=0.265625 nrs=0.140625 sa=7.96719e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=97840 $Y=49910 $D=111
M9058 4095 452 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.1339e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=106810 $Y=35510 $D=111
M9059 VDD 452 4095 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9813e-13 as=1.476e-13 pd=1.89486e-06 ps=1.18e-06 nrd=0.294661 nrs=0.219512 sa=8e-07 sb=6.53902e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=107290 $Y=35510 $D=111
M9060 4094 452 VDD VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.074e-13 as=1.5947e-13 pd=1.96e-06 ps=1.52514e-06 nrd=0.476125 nrs=0.366093 sa=1.24e-06 sb=3.14242e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=107730 $Y=35510 $D=111
M9061 VDD 4094 4096 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.104e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.312909 sa=2.56585e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=108570 $Y=35840 $D=111
M9062 4096 4094 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=7.36585e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=109050 $Y=35840 $D=111
M9063 4097 4098 4096 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.21659e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=109530 $Y=35840 $D=111
M9064 4096 4098 4097 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.69659e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=110010 $Y=35840 $D=111
M9065 4097 418 4095 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.69463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=110950 $Y=35520 $D=111
M9066 4095 418 4097 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=8e-07 sb=1.21463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=111430 $Y=35520 $D=111
M9067 4100 4098 4095 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.28e-06 sb=7.34634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=111910 $Y=35520 $D=111
M9068 4095 4098 4100 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.088e-13 as=1.476e-13 pd=2.36e-06 ps=1.18e-06 nrd=0.310529 nrs=0.219512 sa=1.76e-06 sb=2.54634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=112390 $Y=35520 $D=111
M9069 4100 418 4096 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=3.176e-13 pd=1.18e-06 ps=2.68e-06 nrd=0.219512 nrs=0.472338 sa=3.32683e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=113250 $Y=35840 $D=111
M9070 4096 418 4100 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.4e-13 as=1.476e-13 pd=2.68e-06 ps=1.18e-06 nrd=0.505651 nrs=0.219512 sa=8.12683e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=113730 $Y=35840 $D=111
M9071 VDD 418 4098 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.339e-13 as=3.392e-13 pd=1.69e-06 ps=2.76e-06 nrd=0.29717 nrs=0.301887 sa=3.2e-07 sb=1.91406e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=114790 $Y=35750 $D=111
M9072 4098 418 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.74673e-13 as=3.339e-13 pd=1.84713e-06 ps=1.69e-06 nrd=0.333458 nrs=0.29717 sa=1.07e-06 sb=1.60358e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=115540 $Y=35750 $D=111
M9073 4099 4100 4098 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93608e-13 as=3.39327e-13 pd=1.82905e-06 ps=1.67287e-06 nrd=0.318586 nrs=0.368193 sa=1.86635e-06 sb=1.42469e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=116350 $Y=35860 $D=111
M9074 4102 4097 4099 VDD lppfet w=9.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.20041e-13 as=2.87492e-13 pd=1.66774e-06 ps=1.79095e-06 nrd=0.249028 nrs=0.325364 sa=1.44926e-06 sb=1.38872e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=117010 $Y=35550 $D=111
M9075 4103 4100 4102 VDD lppfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.78404e-13 as=2.15359e-13 pd=1.40371e-06 ps=1.63226e-06 nrd=0.21078 nrs=0.254441 sa=1.4087e-06 sb=1.70522e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=117520 $Y=35890 $D=111
M9076 4101 4097 4103 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.244e-13 as=1.97796e-13 pd=1.46e-06 ps=1.55629e-06 nrd=0.215686 nrs=0.190115 sa=1.39961e-06 sb=1.41e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=118000 $Y=35690 $D=111
M9077 VDD 4102 4101 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.33972e-13 as=2.244e-13 pd=1.57708e-06 ps=1.46e-06 nrd=0.224887 nrs=0.215686 sa=1.6302e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=118560 $Y=35690 $D=111
M9078 4102 446 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.764e-13 as=2.982e-13 pd=3.24e-06 ps=2.01e-06 nrd=0.222722 nrs=0.17645 sa=1.51538e-06 sb=2.89538e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=119120 $Y=35510 $D=111
M9079 VDD 4099 451 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.054e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.247437 sa=3.16719e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=120160 $Y=35510 $D=111
M9080 455 4103 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.352e-13 as=2.304e-13 pd=3.24e-06 ps=1.64e-06 nrd=0.265625 nrs=0.140625 sa=7.96719e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=120640 $Y=35510 $D=111
M9081 4105 413 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.1339e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=110810 $Y=28310 $D=111
M9082 VDD 413 4105 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.9813e-13 as=1.476e-13 pd=1.89486e-06 ps=1.18e-06 nrd=0.294661 nrs=0.219512 sa=8e-07 sb=6.53902e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.44e-14 panw10=0 $X=111290 $Y=28310 $D=111
M9083 4104 413 VDD VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.074e-13 as=1.5947e-13 pd=1.96e-06 ps=1.52514e-06 nrd=0.476125 nrs=0.366093 sa=1.24e-06 sb=3.14242e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=111730 $Y=28310 $D=111
M9084 VDD 4104 4106 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.104e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.312909 sa=2.56585e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=112570 $Y=28640 $D=111
M9085 4106 4104 VDD VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=7.36585e-07 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=113050 $Y=28640 $D=111
M9086 4107 4108 4106 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.21659e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=113530 $Y=28640 $D=111
M9087 4106 4108 4107 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.624e-13 as=1.476e-13 pd=2.28e-06 ps=1.18e-06 nrd=0.390244 nrs=0.219512 sa=1.69659e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=114010 $Y=28640 $D=111
M9088 4107 455 4105 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=2.624e-13 pd=1.18e-06 ps=2.28e-06 nrd=0.219512 nrs=0.390244 sa=3.2e-07 sb=1.69463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=114950 $Y=28320 $D=111
M9089 4105 455 4107 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=8e-07 sb=1.21463e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=115430 $Y=28320 $D=111
M9090 4110 4108 4105 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=1.476e-13 pd=1.18e-06 ps=1.18e-06 nrd=0.219512 nrs=0.219512 sa=1.28e-06 sb=7.34634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=115910 $Y=28320 $D=111
M9091 4105 4108 4110 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.088e-13 as=1.476e-13 pd=2.36e-06 ps=1.18e-06 nrd=0.310529 nrs=0.219512 sa=1.76e-06 sb=2.54634e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=116390 $Y=28320 $D=111
M9092 4110 455 4106 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.476e-13 as=3.176e-13 pd=1.18e-06 ps=2.68e-06 nrd=0.219512 nrs=0.472338 sa=3.32683e-07 sb=8.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=117250 $Y=28640 $D=111
M9093 4106 455 4110 VDD lppfet w=8.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.4e-13 as=1.476e-13 pd=2.68e-06 ps=1.18e-06 nrd=0.505651 nrs=0.219512 sa=8.12683e-07 sb=3.6e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=117730 $Y=28640 $D=111
M9094 VDD 455 4108 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.339e-13 as=3.392e-13 pd=1.69e-06 ps=2.76e-06 nrd=0.29717 nrs=0.301887 sa=3.2e-07 sb=1.91406e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=118790 $Y=28550 $D=111
M9095 4108 455 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.74673e-13 as=3.339e-13 pd=1.84713e-06 ps=1.69e-06 nrd=0.333458 nrs=0.29717 sa=1.07e-06 sb=1.60358e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=7.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=119540 $Y=28550 $D=111
M9096 4109 4110 4108 VDD lppfet w=9.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93608e-13 as=3.39327e-13 pd=1.82905e-06 ps=1.67287e-06 nrd=0.318586 nrs=0.368193 sa=1.86635e-06 sb=1.42469e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=120350 $Y=28660 $D=111
M9097 4112 4107 4109 VDD lppfet w=9.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.20041e-13 as=2.87492e-13 pd=1.66774e-06 ps=1.79095e-06 nrd=0.249028 nrs=0.325364 sa=1.44926e-06 sb=1.38872e-06 sd=0 panw1=0 panw2=1.2e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=121010 $Y=28350 $D=111
M9098 4113 4110 4112 VDD lppfet w=9.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.78404e-13 as=2.15359e-13 pd=1.40371e-06 ps=1.63226e-06 nrd=0.21078 nrs=0.254441 sa=1.4087e-06 sb=1.70522e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=121520 $Y=28690 $D=111
M9099 4111 4107 4113 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.244e-13 as=1.97796e-13 pd=1.46e-06 ps=1.55629e-06 nrd=0.215686 nrs=0.190115 sa=1.39961e-06 sb=1.41e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=122000 $Y=28490 $D=111
M9100 VDD 4112 4111 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.33972e-13 as=2.244e-13 pd=1.57708e-06 ps=1.46e-06 nrd=0.224887 nrs=0.215686 sa=1.6302e-06 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.2e-14 $X=122560 $Y=28490 $D=111
M9101 4112 461 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.764e-13 as=2.982e-13 pd=3.24e-06 ps=2.01e-06 nrd=0.222722 nrs=0.17645 sa=1.51538e-06 sb=2.89538e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=123120 $Y=28310 $D=111
M9102 VDD 4109 463 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.054e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.247437 sa=3.16719e-07 sb=8.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=124160 $Y=28310 $D=111
M9103 448 4113 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.352e-13 as=2.304e-13 pd=3.24e-06 ps=1.64e-06 nrd=0.265625 nrs=0.140625 sa=7.96719e-07 sb=3.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=124640 $Y=28310 $D=111
M9104 4116 30 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3e-13 as=5.2e-13 pd=1.5e-06 ps=3.4e-06 nrd=0.0769231 nrs=0.307692 sa=4e-07 sb=1.58092e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=16940 $Y=49910 $D=111
M9105 4115 43 4116 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.46552e-13 as=1.3e-13 pd=1.86034e-06 ps=1.5e-06 nrd=0.145889 nrs=0.0769231 sa=7.2e-07 sb=1.47262e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=17260 $Y=49910 $D=111
M9106 VDD 61 4115 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92281e-13 as=1.93448e-13 pd=1.49745e-06 ps=1.45966e-06 nrd=0.184814 nrs=0.185936 sa=1.2e-06 sb=1.59529e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.84e-14 panw10=0 $X=17740 $Y=49910 $D=111
M9107 75 4115 VDD VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.892e-13 as=1.62119e-13 pd=1.3e-06 ps=1.26255e-06 nrd=0.255814 nrs=0.219198 sa=1.68e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=18220 $Y=49910 $D=111
M9108 VDD 4115 75 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=1.892e-13 pd=1.22e-06 ps=1.3e-06 nrd=0.209302 nrs=0.255814 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=18780 $Y=49910 $D=111
M9109 75 4115 VDD VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.752e-13 as=1.548e-13 pd=2.36e-06 ps=1.22e-06 nrd=0.372093 nrs=0.209302 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=19260 $Y=49910 $D=111
M9110 4119 431 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.3e-13 as=5.2e-13 pd=1.5e-06 ps=3.4e-06 nrd=0.0769231 nrs=0.307692 sa=4e-07 sb=1.58092e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=109740 $Y=73590 $D=111
M9111 4118 402 4119 VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.46552e-13 as=1.3e-13 pd=1.86034e-06 ps=1.5e-06 nrd=0.145889 nrs=0.0769231 sa=7.2e-07 sb=1.47262e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=110060 $Y=73590 $D=111
M9112 VDD 435 4118 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.92281e-13 as=1.93448e-13 pd=1.49745e-06 ps=1.45966e-06 nrd=0.184814 nrs=0.185936 sa=1.2e-06 sb=1.59529e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.84e-14 panw10=0 $X=110540 $Y=73870 $D=111
M9113 415 4118 VDD VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.892e-13 as=1.62119e-13 pd=1.3e-06 ps=1.26255e-06 nrd=0.255814 nrs=0.219198 sa=1.68e-06 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=111020 $Y=74030 $D=111
M9114 VDD 4118 415 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.548e-13 as=1.892e-13 pd=1.22e-06 ps=1.3e-06 nrd=0.209302 nrs=0.255814 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=111580 $Y=74030 $D=111
M9115 415 4118 VDD VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.752e-13 as=1.548e-13 pd=2.36e-06 ps=1.22e-06 nrd=0.372093 nrs=0.209302 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.92e-14 panw10=0 $X=112060 $Y=74030 $D=111
M9116 4121 74 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=3.549e-13 pd=1.04e-06 ps=2.715e-06 nrd=0.119048 nrs=0.502976 sa=3.6e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=23790 $Y=28430 $D=111
M9117 77 57 4121 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=24110 $Y=28430 $D=111
M9118 4122 84 77 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.16e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=24590 $Y=28430 $D=111
M9119 VDD 83 4122 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.801e-13 as=8.4e-14 pd=2.775e-06 ps=1.04e-06 nrd=0.53869 nrs=0.119048 sa=1.48e-06 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=24910 $Y=28430 $D=111
M9120 4124 102 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=3.549e-13 pd=1.04e-06 ps=2.715e-06 nrd=0.119048 nrs=0.502976 sa=3.6e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=29790 $Y=30730 $D=111
M9121 106 74 4124 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=30110 $Y=30730 $D=111
M9122 4125 84 106 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.16e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=30590 $Y=30730 $D=111
M9123 VDD 112 4125 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.801e-13 as=8.4e-14 pd=2.775e-06 ps=1.04e-06 nrd=0.53869 nrs=0.119048 sa=1.48e-06 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=30910 $Y=30730 $D=111
M9124 4127 148 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=3.549e-13 pd=1.04e-06 ps=2.715e-06 nrd=0.119048 nrs=0.502976 sa=3.6e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=38590 $Y=23530 $D=111
M9125 155 144 4127 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=38910 $Y=23530 $D=111
M9126 4128 182 155 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.16e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=39390 $Y=23530 $D=111
M9127 VDD 165 4128 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.801e-13 as=8.4e-14 pd=2.775e-06 ps=1.04e-06 nrd=0.53869 nrs=0.119048 sa=1.48e-06 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=39710 $Y=23530 $D=111
M9128 4130 148 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=3.549e-13 pd=1.04e-06 ps=2.715e-06 nrd=0.119048 nrs=0.502976 sa=3.6e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=40190 $Y=50030 $D=111
M9129 178 166 4130 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=40510 $Y=50030 $D=111
M9130 4131 164 178 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.16e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=40990 $Y=50030 $D=111
M9131 VDD 198 4131 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.801e-13 as=8.4e-14 pd=2.775e-06 ps=1.04e-06 nrd=0.53869 nrs=0.119048 sa=1.48e-06 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=41310 $Y=50030 $D=111
M9132 4133 148 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=3.549e-13 pd=1.04e-06 ps=2.715e-06 nrd=0.119048 nrs=0.502976 sa=3.6e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=42590 $Y=35630 $D=111
M9133 93 164 4133 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=42910 $Y=35630 $D=111
M9134 4134 198 93 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.16e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=43390 $Y=35630 $D=111
M9135 VDD 144 4134 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.801e-13 as=8.4e-14 pd=2.775e-06 ps=1.04e-06 nrd=0.53869 nrs=0.119048 sa=1.48e-06 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=43710 $Y=35630 $D=111
M9136 4136 293 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=3.549e-13 pd=1.04e-06 ps=2.715e-06 nrd=0.119048 nrs=0.502976 sa=3.6e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=73390 $Y=57230 $D=111
M9137 288 325 4136 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=73710 $Y=57230 $D=111
M9138 4137 295 288 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.16e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=74190 $Y=57230 $D=111
M9139 VDD 280 4137 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.801e-13 as=8.4e-14 pd=2.775e-06 ps=1.04e-06 nrd=0.53869 nrs=0.119048 sa=1.48e-06 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=74510 $Y=57230 $D=111
M9140 4139 343 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=3.549e-13 pd=1.04e-06 ps=2.715e-06 nrd=0.119048 nrs=0.502976 sa=3.6e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=88590 $Y=52330 $D=111
M9141 331 325 4139 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=88910 $Y=52330 $D=111
M9142 4140 295 331 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.16e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=89390 $Y=52330 $D=111
M9143 VDD 328 4140 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.801e-13 as=8.4e-14 pd=2.775e-06 ps=1.04e-06 nrd=0.53869 nrs=0.119048 sa=1.48e-06 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=89710 $Y=52330 $D=111
M9144 4142 400 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=3.549e-13 pd=1.04e-06 ps=2.715e-06 nrd=0.119048 nrs=0.502976 sa=3.6e-07 sb=1.52e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=108190 $Y=45130 $D=111
M9145 910 406 4142 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.512e-13 as=8.4e-14 pd=1.2e-06 ps=1.04e-06 nrd=0.214286 nrs=0.119048 sa=6.8e-07 sb=1.2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=108510 $Y=45130 $D=111
M9146 4143 416 910 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=8.4e-14 as=1.512e-13 pd=1.04e-06 ps=1.2e-06 nrd=0.119048 nrs=0.214286 sa=1.16e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=108990 $Y=45130 $D=111
M9147 VDD 410 4143 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.801e-13 as=8.4e-14 pd=2.775e-06 ps=1.04e-06 nrd=0.53869 nrs=0.119048 sa=1.48e-06 sb=4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=3.6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.12e-14 panw10=0 $X=109310 $Y=45130 $D=111
M9148 4145 84 70 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=17640 $Y=35690 $D=111
M9149 VDD 57 4145 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=17960 $Y=35690 $D=111
M9150 4146 57 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=18440 $Y=35690 $D=111
M9151 70 84 4146 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=18760 $Y=35690 $D=111
M9152 4147 84 70 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=19240 $Y=35690 $D=111
M9153 VDD 57 4147 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=19560 $Y=35690 $D=111
M9154 4148 142 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=20040 $Y=35690 $D=111
M9155 70 74 4148 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=20360 $Y=35690 $D=111
M9156 4149 74 70 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=20840 $Y=35690 $D=111
M9157 VDD 142 4149 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=21160 $Y=35690 $D=111
M9158 4150 142 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=21640 $Y=35690 $D=111
M9159 70 74 4150 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=21960 $Y=35690 $D=111
M9160 4152 181 273 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=44840 $Y=59190 $D=111
M9161 VDD 189 4152 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=45160 $Y=59190 $D=111
M9162 4153 189 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=45640 $Y=59190 $D=111
M9163 273 181 4153 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=45960 $Y=59190 $D=111
M9164 4154 181 273 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=46440 $Y=59190 $D=111
M9165 VDD 189 4154 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=46760 $Y=59190 $D=111
M9166 4155 179 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=47240 $Y=59190 $D=111
M9167 273 151 4155 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=47560 $Y=59190 $D=111
M9168 4156 151 273 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=48040 $Y=59190 $D=111
M9169 VDD 179 4156 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=48360 $Y=59190 $D=111
M9170 4157 179 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=48840 $Y=59190 $D=111
M9171 273 151 4157 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=49160 $Y=59190 $D=111
M9172 4159 212 194 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=52840 $Y=37590 $D=111
M9173 VDD 199 4159 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=53160 $Y=37590 $D=111
M9174 4160 199 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=53640 $Y=37590 $D=111
M9175 194 212 4160 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=53960 $Y=37590 $D=111
M9176 4161 212 194 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=54440 $Y=37590 $D=111
M9177 VDD 199 4161 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=54760 $Y=37590 $D=111
M9178 4162 219 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=55240 $Y=37590 $D=111
M9179 194 232 4162 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=55560 $Y=37590 $D=111
M9180 4163 232 194 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=56040 $Y=37590 $D=111
M9181 VDD 219 4163 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=56360 $Y=37590 $D=111
M9182 4164 219 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=56840 $Y=37590 $D=111
M9183 194 232 4164 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=57160 $Y=37590 $D=111
M9184 4166 199 224 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=61240 $Y=35690 $D=111
M9185 VDD 209 4166 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=61560 $Y=35690 $D=111
M9186 4167 209 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=62040 $Y=35690 $D=111
M9187 224 199 4167 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=62360 $Y=35690 $D=111
M9188 4168 199 224 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=62840 $Y=35690 $D=111
M9189 VDD 209 4168 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=63160 $Y=35690 $D=111
M9190 4169 231 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=63640 $Y=35690 $D=111
M9191 224 242 4169 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=63960 $Y=35690 $D=111
M9192 4170 242 224 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=64440 $Y=35690 $D=111
M9193 VDD 231 4170 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=64760 $Y=35690 $D=111
M9194 4171 231 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=65240 $Y=35690 $D=111
M9195 224 242 4171 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=65560 $Y=35690 $D=111
M9196 4173 301 279 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=69640 $Y=37590 $D=111
M9197 VDD 267 4173 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=69960 $Y=37590 $D=111
M9198 4174 267 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=70440 $Y=37590 $D=111
M9199 279 301 4174 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=70760 $Y=37590 $D=111
M9200 4175 301 279 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=71240 $Y=37590 $D=111
M9201 VDD 267 4175 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=71560 $Y=37590 $D=111
M9202 4176 212 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=72040 $Y=37590 $D=111
M9203 279 282 4176 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=72360 $Y=37590 $D=111
M9204 4177 282 279 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=72840 $Y=37590 $D=111
M9205 VDD 212 4177 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=73160 $Y=37590 $D=111
M9206 4178 212 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=73640 $Y=37590 $D=111
M9207 279 282 4178 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=73960 $Y=37590 $D=111
M9208 4180 328 341 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=74840 $Y=50090 $D=111
M9209 VDD 325 4180 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=75160 $Y=50090 $D=111
M9210 4181 325 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=75640 $Y=50090 $D=111
M9211 341 328 4181 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=75960 $Y=50090 $D=111
M9212 4182 328 341 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=76440 $Y=50090 $D=111
M9213 VDD 325 4182 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=76760 $Y=50090 $D=111
M9214 4183 293 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=77240 $Y=50090 $D=111
M9215 341 295 4183 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=77560 $Y=50090 $D=111
M9216 4184 295 341 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=78040 $Y=50090 $D=111
M9217 VDD 293 4184 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=78360 $Y=50090 $D=111
M9218 4185 293 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=78840 $Y=50090 $D=111
M9219 341 295 4185 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=79160 $Y=50090 $D=111
M9220 4187 314 346 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=89640 $Y=35690 $D=111
M9221 VDD 336 4187 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=89960 $Y=35690 $D=111
M9222 4188 336 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=90440 $Y=35690 $D=111
M9223 346 314 4188 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=90760 $Y=35690 $D=111
M9224 4189 314 346 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=91240 $Y=35690 $D=111
M9225 VDD 336 4189 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=91560 $Y=35690 $D=111
M9226 4190 327 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=92040 $Y=35690 $D=111
M9227 346 330 4190 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=92360 $Y=35690 $D=111
M9228 4191 330 346 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=92840 $Y=35690 $D=111
M9229 VDD 327 4191 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=93160 $Y=35690 $D=111
M9230 4192 327 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=93640 $Y=35690 $D=111
M9231 346 330 4192 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=93960 $Y=35690 $D=111
M9232 4194 336 348 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=92040 $Y=42890 $D=111
M9233 VDD 327 4194 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=92360 $Y=42890 $D=111
M9234 4195 327 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=92840 $Y=42890 $D=111
M9235 348 336 4195 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=93160 $Y=42890 $D=111
M9236 4196 336 348 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=93640 $Y=42890 $D=111
M9237 VDD 327 4196 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=93960 $Y=42890 $D=111
M9238 4197 319 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=94440 $Y=42890 $D=111
M9239 348 330 4197 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=94760 $Y=42890 $D=111
M9240 4198 330 348 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=95240 $Y=42890 $D=111
M9241 VDD 319 4198 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=95560 $Y=42890 $D=111
M9242 4199 319 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=96040 $Y=42890 $D=111
M9243 348 330 4199 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=96360 $Y=42890 $D=111
M9244 4201 419 365 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=3.584e-13 pd=1.32e-06 ps=2.88e-06 nrd=0.0892857 nrs=0.285714 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=108040 $Y=42890 $D=111
M9245 VDD 400 4201 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=6.4e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=108360 $Y=42890 $D=111
M9246 4202 400 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.12e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=108840 $Y=42890 $D=111
M9247 365 419 4202 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=1.44e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=109160 $Y=42890 $D=111
M9248 4203 419 365 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=1.92e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=109640 $Y=42890 $D=111
M9249 VDD 400 4203 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=109960 $Y=42890 $D=111
M9250 4204 343 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=110440 $Y=42890 $D=111
M9251 365 410 4204 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.92e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=110760 $Y=42890 $D=111
M9252 4205 410 365 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=1.44e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=111240 $Y=42890 $D=111
M9253 VDD 343 4205 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.016e-13 as=1.12e-13 pd=1.48e-06 ps=1.32e-06 nrd=0.160714 nrs=0.0892857 sa=2e-06 sb=1.12e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=111560 $Y=42890 $D=111
M9254 4206 343 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12e-13 as=2.016e-13 pd=1.32e-06 ps=1.48e-06 nrd=0.0892857 nrs=0.160714 sa=2e-06 sb=6.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=112040 $Y=42890 $D=111
M9255 365 410 4206 VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.584e-13 as=1.12e-13 pd=2.88e-06 ps=1.32e-06 nrd=0.285714 nrs=0.0892857 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=2.4e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=112360 $Y=42890 $D=111
M9256 VDD 148 4207 VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26104e-13 as=2.176e-13 pd=1.10627e-06 ps=2e-06 nrd=0.272717 nrs=0.470588 sa=3.2e-07 sb=1.17603e-06 sd=0 panw1=0 panw2=4.5e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.22e-14 panw9=9e-16 panw10=0 $X=53450 $Y=57110 $D=111
M9257 VDD 4208 234 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.944e-13 pd=1.6e-06 ps=3.2e-06 nrd=0.125 nrs=0.179687 sa=2.3e-07 sb=9.59531e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=1.536e-13 $X=53650 $Y=58240 $D=111
M9258 4207 168 VDD VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=1.22396e-13 pd=1.02e-06 ps=1.07373e-06 nrd=0.272727 nrs=0.280981 sa=7.54545e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=53930 $Y=57060 $D=111
M9259 4208 200 4207 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.112e-13 as=1.188e-13 pd=1.96e-06 ps=1.02e-06 nrd=0.484848 nrs=0.272727 sa=1.23455e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=54410 $Y=57060 $D=111
M9260 VDD 400 4210 VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.26104e-13 as=2.176e-13 pd=1.10627e-06 ps=2e-06 nrd=0.272717 nrs=0.470588 sa=3.2e-07 sb=1.17603e-06 sd=0 panw1=0 panw2=4.5e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.22e-14 panw9=9e-16 panw10=0 $X=105450 $Y=45410 $D=111
M9261 403 4211 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.944e-13 as=2.048e-13 pd=3.2e-06 ps=1.6e-06 nrd=0.179687 nrs=0.125 sa=7.41328e-07 sb=2.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=1.536e-13 $X=105650 $Y=44840 $D=111
M9262 4210 410 VDD VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.188e-13 as=1.22396e-13 pd=1.02e-06 ps=1.07373e-06 nrd=0.272727 nrs=0.280981 sa=7.54545e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=105930 $Y=45480 $D=111
M9263 4211 406 4210 VDD lppfet w=6.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.112e-13 as=1.188e-13 pd=1.96e-06 ps=1.02e-06 nrd=0.484848 nrs=0.272727 sa=1.23455e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.92e-14 panw9=0 panw10=0 $X=106410 $Y=45480 $D=111
M9264 110 89 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=4.064e-13 pd=1.63e-06 ps=3.18e-06 nrd=0.141732 nrs=0.251969 sa=3.2e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.04e-14 $X=32900 $Y=64310 $D=111
M9265 VDD 89 110 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.38846e-13 as=2.286e-13 pd=3.12994e-06 ps=1.63e-06 nrd=0.272085 nrs=0.141732 sa=8e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.04e-14 $X=33380 $Y=64310 $D=111
M9266 371 344 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=4.064e-13 pd=1.63e-06 ps=3.18e-06 nrd=0.141732 nrs=0.251969 sa=3.2e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.04e-14 $X=100900 $Y=13910 $D=111
M9267 VDD 344 371 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.38846e-13 as=2.286e-13 pd=3.12994e-06 ps=1.63e-06 nrd=0.272085 nrs=0.141732 sa=8e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.04e-14 $X=101380 $Y=13910 $D=111
M9268 VDD 150 4215 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.69778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=7.8e-14 panw8=9.96e-14 panw9=4.56e-14 panw10=0 $X=8810 $Y=45010 $D=111
M9269 4215 150 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.21778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.752e-13 panw10=0 $X=9290 $Y=45010 $D=111
M9270 VDD 150 4215 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.96397e-13 as=1.944e-13 pd=1.50655e-06 ps=1.44e-06 nrd=0.168378 nrs=0.166667 sa=1.28e-06 sb=7.37778e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=1.296e-13 $X=9770 $Y=45010 $D=111
M9271 4213 150 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.36403e-13 pd=3.24e-06 ps=1.81345e-06 nrd=0.190769 nrs=0.139884 sa=1.496e-06 sb=2.48e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=10250 $Y=44790 $D=111
M9272 4216 4213 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=2.496e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.213992 sa=2.31111e-07 sb=1.73556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=11070 $Y=45110 $D=111
M9273 VDD 4213 4216 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=7.11111e-07 sb=1.58444e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=11550 $Y=45110 $D=111
M9274 4216 4213 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.12366e-13 as=1.944e-13 pd=1.77645e-06 ps=1.44e-06 nrd=0.18207 nrs=0.166667 sa=1.19111e-06 sb=1.43333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=12030 $Y=45110 $D=111
M9275 4217 4214 4216 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.08434e-13 pd=1.42e-06 ps=1.74355e-06 nrd=0.169811 nrs=0.185505 sa=1.25811e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=2e-15 panw7=2.08e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3.24e-14 $X=12510 $Y=44790 $D=111
M9276 4216 4214 4217 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.62264e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=12990 $Y=44790 $D=111
M9277 4217 4214 4216 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.76755e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=13470 $Y=44790 $D=111
M9278 4215 53 4217 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.91245e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=13950 $Y=44790 $D=111
M9279 4217 53 4215 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=14430 $Y=44790 $D=111
M9280 4215 53 4217 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=14910 $Y=44790 $D=111
M9281 4218 4214 4215 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=15390 $Y=44790 $D=111
M9282 4215 4214 4218 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.738e-13 as=1.908e-13 pd=1.79e-06 ps=1.42e-06 nrd=0.243681 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=15870 $Y=44790 $D=111
M9283 4218 4214 4215 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.738e-13 pd=1.42e-06 ps=1.79e-06 nrd=0.169811 nrs=0.243681 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=16430 $Y=44790 $D=111
M9284 4216 53 4218 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=16910 $Y=44790 $D=111
M9285 4218 53 4216 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=17390 $Y=44790 $D=111
M9286 4216 53 4218 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=1.908e-13 pd=2.76e-06 ps=1.42e-06 nrd=0.301887 nrs=0.169811 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=17870 $Y=44790 $D=111
M9287 VDD 53 4214 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.96111e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=18990 $Y=44790 $D=111
M9288 4214 53 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.89444e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=19470 $Y=44790 $D=111
M9289 VDD 53 4214 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=1.28e-06 sb=1.60574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=19950 $Y=44790 $D=111
M9290 4214 53 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.0246e-13 as=1.944e-13 pd=1.54746e-06 ps=1.44e-06 nrd=0.173577 nrs=0.166667 sa=1.76e-06 sb=1.12574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=20430 $Y=44790 $D=111
M9291 4219 4218 4214 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.7434e-13 pd=1.29e-06 ps=1.33254e-06 nrd=0.193548 nrs=0.201573 sa=2e-06 sb=7.82151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=20910 $Y=44940 $D=111
M9292 4214 4218 4219 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.81e-13 as=1.674e-13 pd=2.66e-06 ps=1.29e-06 nrd=0.324893 nrs=0.193548 sa=2e-06 sb=3.02151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=21390 $Y=44940 $D=111
M9293 4221 4217 4219 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.756e-13 pd=9.8e-07 ps=1.96e-06 nrd=0.290323 nrs=0.456816 sa=2.83226e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=22310 $Y=45110 $D=111
M9294 4219 4217 4221 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.116e-13 pd=9.8e-07 ps=9.8e-07 nrd=0.290323 nrs=0.290323 sa=7.63226e-07 sb=1.79742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=22790 $Y=45110 $D=111
M9295 4221 4217 4219 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24e-13 as=1.116e-13 pd=1.032e-06 ps=9.8e-07 nrd=0.322581 nrs=0.290323 sa=1.24323e-06 sb=1.31742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=23270 $Y=45110 $D=111
M9296 4222 4218 4221 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.86e-13 pd=1.29e-06 ps=1.548e-06 nrd=0.193548 nrs=0.215054 sa=1.24215e-06 sb=7.84946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=23750 $Y=44800 $D=111
M9297 4221 4218 4222 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.424e-13 as=1.674e-13 pd=3e-06 ps=1.29e-06 nrd=0.395884 nrs=0.193548 sa=1.58667e-06 sb=3.04946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=24230 $Y=44800 $D=111
M9298 4222 4217 4220 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=2.844e-13 pd=1.29e-06 ps=2.5e-06 nrd=0.193548 nrs=0.328824 sa=3.05806e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=25440 $Y=45010 $D=111
M9299 4220 4217 4222 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.674e-13 pd=1.29e-06 ps=1.29e-06 nrd=0.193548 nrs=0.193548 sa=7.85806e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=25920 $Y=45010 $D=111
M9300 VDD 4221 4220 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30175e-13 as=1.674e-13 pd=1.54446e-06 ps=1.29e-06 nrd=0.266129 nrs=0.193548 sa=1.26581e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=26400 $Y=45010 $D=111
M9301 4220 4221 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.296e-13 as=2.54925e-13 pd=2.7e-06 ps=1.71054e-06 nrd=0.31068 nrs=0.240291 sa=1.6835e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=26960 $Y=44910 $D=111
M9302 VDD 94 4221 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.90115e-13 as=4.128e-13 pd=1.8042e-06 ps=3.22e-06 nrd=0.174337 nrs=0.248062 sa=3.2e-07 sb=8.34419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=27900 $Y=44790 $D=111
M9303 4221 94 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.54e-13 as=2.90115e-13 pd=3.22e-06 ps=1.8042e-06 nrd=0.212728 nrs=0.174337 sa=8.8e-07 sb=2.74419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=28460 $Y=44790 $D=111
M9304 44 4219 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=29560 $Y=44800 $D=111
M9305 VDD 4219 44 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=30040 $Y=44800 $D=111
M9306 21 4222 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.56e-13 as=2.304e-13 pd=1.68e-06 ps=1.64e-06 nrd=0.15625 nrs=0.140625 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=30520 $Y=44800 $D=111
M9307 VDD 4222 21 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.56e-13 pd=3.2e-06 ps=1.68e-06 nrd=0.25 nrs=0.15625 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=31040 $Y=44800 $D=111
M9308 VDD 103 4225 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.69778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=28010 $Y=37810 $D=111
M9309 4225 103 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.21778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=28490 $Y=37810 $D=111
M9310 VDD 103 4225 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.96397e-13 as=1.944e-13 pd=1.50655e-06 ps=1.44e-06 nrd=0.168378 nrs=0.166667 sa=1.28e-06 sb=7.37778e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=28970 $Y=37810 $D=111
M9311 4223 103 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.36403e-13 pd=3.24e-06 ps=1.81345e-06 nrd=0.190769 nrs=0.139884 sa=1.496e-06 sb=2.48e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=29450 $Y=37590 $D=111
M9312 4226 4223 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=2.496e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.213992 sa=2.31111e-07 sb=1.73556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=30270 $Y=37910 $D=111
M9313 VDD 4223 4226 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=7.11111e-07 sb=1.58444e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=30750 $Y=37910 $D=111
M9314 4226 4223 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.12366e-13 as=1.944e-13 pd=1.77645e-06 ps=1.44e-06 nrd=0.18207 nrs=0.166667 sa=1.19111e-06 sb=1.43333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=31230 $Y=37910 $D=111
M9315 4227 4224 4226 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.08434e-13 pd=1.42e-06 ps=1.74355e-06 nrd=0.169811 nrs=0.185505 sa=1.25811e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=2e-15 panw7=2.08e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3.24e-14 $X=31710 $Y=37590 $D=111
M9316 4226 4224 4227 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.62264e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=32190 $Y=37590 $D=111
M9317 4227 4224 4226 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.76755e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=32670 $Y=37590 $D=111
M9318 4225 194 4227 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.91245e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=33150 $Y=37590 $D=111
M9319 4227 194 4225 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=33630 $Y=37590 $D=111
M9320 4225 194 4227 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=34110 $Y=37590 $D=111
M9321 4228 4224 4225 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=34590 $Y=37590 $D=111
M9322 4225 4224 4228 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.738e-13 as=1.908e-13 pd=1.79e-06 ps=1.42e-06 nrd=0.243681 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=35070 $Y=37590 $D=111
M9323 4228 4224 4225 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.738e-13 pd=1.42e-06 ps=1.79e-06 nrd=0.169811 nrs=0.243681 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=35630 $Y=37590 $D=111
M9324 4226 194 4228 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=36110 $Y=37590 $D=111
M9325 4228 194 4226 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=36590 $Y=37590 $D=111
M9326 4226 194 4228 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=1.908e-13 pd=2.76e-06 ps=1.42e-06 nrd=0.301887 nrs=0.169811 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=37070 $Y=37590 $D=111
M9327 VDD 194 4224 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.96111e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=38190 $Y=37590 $D=111
M9328 4224 194 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.89444e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=38670 $Y=37590 $D=111
M9329 VDD 194 4224 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=1.28e-06 sb=1.60574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=39150 $Y=37590 $D=111
M9330 4224 194 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.0246e-13 as=1.944e-13 pd=1.54746e-06 ps=1.44e-06 nrd=0.173577 nrs=0.166667 sa=1.76e-06 sb=1.12574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=39630 $Y=37590 $D=111
M9331 4229 4228 4224 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.7434e-13 pd=1.29e-06 ps=1.33254e-06 nrd=0.193548 nrs=0.201573 sa=2e-06 sb=7.82151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=40110 $Y=37740 $D=111
M9332 4224 4228 4229 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.81e-13 as=1.674e-13 pd=2.66e-06 ps=1.29e-06 nrd=0.324893 nrs=0.193548 sa=2e-06 sb=3.02151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=40590 $Y=37740 $D=111
M9333 4231 4227 4229 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.756e-13 pd=9.8e-07 ps=1.96e-06 nrd=0.290323 nrs=0.456816 sa=2.83226e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=41510 $Y=37910 $D=111
M9334 4229 4227 4231 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.116e-13 pd=9.8e-07 ps=9.8e-07 nrd=0.290323 nrs=0.290323 sa=7.63226e-07 sb=1.79742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=41990 $Y=37910 $D=111
M9335 4231 4227 4229 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24e-13 as=1.116e-13 pd=1.032e-06 ps=9.8e-07 nrd=0.322581 nrs=0.290323 sa=1.24323e-06 sb=1.31742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=42470 $Y=37910 $D=111
M9336 4232 4228 4231 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.86e-13 pd=1.29e-06 ps=1.548e-06 nrd=0.193548 nrs=0.215054 sa=1.24215e-06 sb=7.84946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=42950 $Y=37600 $D=111
M9337 4231 4228 4232 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.424e-13 as=1.674e-13 pd=3e-06 ps=1.29e-06 nrd=0.395884 nrs=0.193548 sa=1.58667e-06 sb=3.04946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=43430 $Y=37600 $D=111
M9338 4232 4227 4230 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=2.844e-13 pd=1.29e-06 ps=2.5e-06 nrd=0.193548 nrs=0.328824 sa=3.05806e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=44640 $Y=37810 $D=111
M9339 4230 4227 4232 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.674e-13 pd=1.29e-06 ps=1.29e-06 nrd=0.193548 nrs=0.193548 sa=7.85806e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=45120 $Y=37810 $D=111
M9340 VDD 4231 4230 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30175e-13 as=1.674e-13 pd=1.54446e-06 ps=1.29e-06 nrd=0.266129 nrs=0.193548 sa=1.26581e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=45600 $Y=37810 $D=111
M9341 4230 4231 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.296e-13 as=2.54925e-13 pd=2.7e-06 ps=1.71054e-06 nrd=0.31068 nrs=0.240291 sa=1.6835e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=46160 $Y=37710 $D=111
M9342 VDD 178 4231 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.90115e-13 as=4.128e-13 pd=1.8042e-06 ps=3.22e-06 nrd=0.174337 nrs=0.248062 sa=3.2e-07 sb=8.34419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=47100 $Y=37590 $D=111
M9343 4231 178 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.54e-13 as=2.90115e-13 pd=3.22e-06 ps=1.8042e-06 nrd=0.212728 nrs=0.174337 sa=8.8e-07 sb=2.74419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=47660 $Y=37590 $D=111
M9344 120 4229 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=48760 $Y=37600 $D=111
M9345 VDD 4229 120 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=49240 $Y=37600 $D=111
M9346 94 4232 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.56e-13 as=2.304e-13 pd=1.68e-06 ps=1.64e-06 nrd=0.15625 nrs=0.140625 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=49720 $Y=37600 $D=111
M9347 VDD 4232 94 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.56e-13 pd=3.2e-06 ps=1.68e-06 nrd=0.25 nrs=0.15625 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=50240 $Y=37600 $D=111
M9348 VDD 253 4235 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.69778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=54010 $Y=66610 $D=111
M9349 4235 253 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.21778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=54490 $Y=66610 $D=111
M9350 VDD 253 4235 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.96397e-13 as=1.944e-13 pd=1.50655e-06 ps=1.44e-06 nrd=0.168378 nrs=0.166667 sa=1.28e-06 sb=7.37778e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=54970 $Y=66610 $D=111
M9351 4233 253 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.36403e-13 pd=3.24e-06 ps=1.81345e-06 nrd=0.190769 nrs=0.139884 sa=1.496e-06 sb=2.48e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=55450 $Y=66390 $D=111
M9352 4236 4233 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=2.496e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.213992 sa=2.31111e-07 sb=1.73556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=56270 $Y=66710 $D=111
M9353 VDD 4233 4236 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=7.11111e-07 sb=1.58444e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=56750 $Y=66710 $D=111
M9354 4236 4233 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.12366e-13 as=1.944e-13 pd=1.77645e-06 ps=1.44e-06 nrd=0.18207 nrs=0.166667 sa=1.19111e-06 sb=1.43333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=57230 $Y=66710 $D=111
M9355 4237 4234 4236 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.08434e-13 pd=1.42e-06 ps=1.74355e-06 nrd=0.169811 nrs=0.185505 sa=1.25811e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=2e-15 panw7=2.08e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3.24e-14 $X=57710 $Y=66390 $D=111
M9356 4236 4234 4237 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.62264e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=58190 $Y=66390 $D=111
M9357 4237 4234 4236 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.76755e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=58670 $Y=66390 $D=111
M9358 4235 276 4237 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.91245e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=59150 $Y=66390 $D=111
M9359 4237 276 4235 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=59630 $Y=66390 $D=111
M9360 4235 276 4237 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=60110 $Y=66390 $D=111
M9361 4238 4234 4235 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=60590 $Y=66390 $D=111
M9362 4235 4234 4238 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.738e-13 as=1.908e-13 pd=1.79e-06 ps=1.42e-06 nrd=0.243681 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=61070 $Y=66390 $D=111
M9363 4238 4234 4235 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.738e-13 pd=1.42e-06 ps=1.79e-06 nrd=0.169811 nrs=0.243681 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=61630 $Y=66390 $D=111
M9364 4236 276 4238 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=62110 $Y=66390 $D=111
M9365 4238 276 4236 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=62590 $Y=66390 $D=111
M9366 4236 276 4238 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=1.908e-13 pd=2.76e-06 ps=1.42e-06 nrd=0.301887 nrs=0.169811 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=63070 $Y=66390 $D=111
M9367 VDD 276 4234 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.96111e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=64190 $Y=66390 $D=111
M9368 4234 276 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.89444e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=64670 $Y=66390 $D=111
M9369 VDD 276 4234 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=1.28e-06 sb=1.60574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=65150 $Y=66390 $D=111
M9370 4234 276 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.0246e-13 as=1.944e-13 pd=1.54746e-06 ps=1.44e-06 nrd=0.173577 nrs=0.166667 sa=1.76e-06 sb=1.12574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=65630 $Y=66390 $D=111
M9371 4239 4238 4234 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.7434e-13 pd=1.29e-06 ps=1.33254e-06 nrd=0.193548 nrs=0.201573 sa=2e-06 sb=7.82151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=66110 $Y=66540 $D=111
M9372 4234 4238 4239 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.81e-13 as=1.674e-13 pd=2.66e-06 ps=1.29e-06 nrd=0.324893 nrs=0.193548 sa=2e-06 sb=3.02151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=66590 $Y=66540 $D=111
M9373 4241 4237 4239 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.756e-13 pd=9.8e-07 ps=1.96e-06 nrd=0.290323 nrs=0.456816 sa=2.83226e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=67510 $Y=66710 $D=111
M9374 4239 4237 4241 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.116e-13 pd=9.8e-07 ps=9.8e-07 nrd=0.290323 nrs=0.290323 sa=7.63226e-07 sb=1.79742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=67990 $Y=66710 $D=111
M9375 4241 4237 4239 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24e-13 as=1.116e-13 pd=1.032e-06 ps=9.8e-07 nrd=0.322581 nrs=0.290323 sa=1.24323e-06 sb=1.31742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=68470 $Y=66710 $D=111
M9376 4242 4238 4241 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.86e-13 pd=1.29e-06 ps=1.548e-06 nrd=0.193548 nrs=0.215054 sa=1.24215e-06 sb=7.84946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=68950 $Y=66400 $D=111
M9377 4241 4238 4242 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.424e-13 as=1.674e-13 pd=3e-06 ps=1.29e-06 nrd=0.395884 nrs=0.193548 sa=1.58667e-06 sb=3.04946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=69430 $Y=66400 $D=111
M9378 4242 4237 4240 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=2.844e-13 pd=1.29e-06 ps=2.5e-06 nrd=0.193548 nrs=0.328824 sa=3.05806e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=70640 $Y=66610 $D=111
M9379 4240 4237 4242 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.674e-13 pd=1.29e-06 ps=1.29e-06 nrd=0.193548 nrs=0.193548 sa=7.85806e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=71120 $Y=66610 $D=111
M9380 VDD 4241 4240 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30175e-13 as=1.674e-13 pd=1.54446e-06 ps=1.29e-06 nrd=0.266129 nrs=0.193548 sa=1.26581e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=71600 $Y=66610 $D=111
M9381 4240 4241 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.296e-13 as=2.54925e-13 pd=2.7e-06 ps=1.71054e-06 nrd=0.31068 nrs=0.240291 sa=1.6835e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=72160 $Y=66510 $D=111
M9382 VDD 275 4241 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.90115e-13 as=4.128e-13 pd=1.8042e-06 ps=3.22e-06 nrd=0.174337 nrs=0.248062 sa=3.2e-07 sb=8.34419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=73100 $Y=66390 $D=111
M9383 4241 275 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.54e-13 as=2.90115e-13 pd=3.22e-06 ps=1.8042e-06 nrd=0.212728 nrs=0.174337 sa=8.8e-07 sb=2.74419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=73660 $Y=66390 $D=111
M9384 309 4239 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=74760 $Y=66400 $D=111
M9385 VDD 4239 309 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=75240 $Y=66400 $D=111
M9386 289 4242 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.56e-13 as=2.304e-13 pd=1.68e-06 ps=1.64e-06 nrd=0.15625 nrs=0.140625 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=75720 $Y=66400 $D=111
M9387 VDD 4242 289 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.56e-13 pd=3.2e-06 ps=1.68e-06 nrd=0.25 nrs=0.15625 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=76240 $Y=66400 $D=111
M9388 VDD 234 4245 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.69778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=63610 $Y=52210 $D=111
M9389 4245 234 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.21778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=64090 $Y=52210 $D=111
M9390 VDD 234 4245 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.96397e-13 as=1.944e-13 pd=1.50655e-06 ps=1.44e-06 nrd=0.168378 nrs=0.166667 sa=1.28e-06 sb=7.37778e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=64570 $Y=52210 $D=111
M9391 4243 234 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.36403e-13 pd=3.24e-06 ps=1.81345e-06 nrd=0.190769 nrs=0.139884 sa=1.496e-06 sb=2.48e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=65050 $Y=51990 $D=111
M9392 4246 4243 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=2.496e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.213992 sa=2.31111e-07 sb=1.73556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=65870 $Y=52310 $D=111
M9393 VDD 4243 4246 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=7.11111e-07 sb=1.58444e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=66350 $Y=52310 $D=111
M9394 4246 4243 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.12366e-13 as=1.944e-13 pd=1.77645e-06 ps=1.44e-06 nrd=0.18207 nrs=0.166667 sa=1.19111e-06 sb=1.43333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=66830 $Y=52310 $D=111
M9395 4247 4244 4246 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.08434e-13 pd=1.42e-06 ps=1.74355e-06 nrd=0.169811 nrs=0.185505 sa=1.25811e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=2e-15 panw7=2.08e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3.24e-14 $X=67310 $Y=51990 $D=111
M9396 4246 4244 4247 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.62264e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=67790 $Y=51990 $D=111
M9397 4247 4244 4246 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.76755e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=68270 $Y=51990 $D=111
M9398 4245 824 4247 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.91245e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=68750 $Y=51990 $D=111
M9399 4247 824 4245 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=69230 $Y=51990 $D=111
M9400 4245 824 4247 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=69710 $Y=51990 $D=111
M9401 4248 4244 4245 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=70190 $Y=51990 $D=111
M9402 4245 4244 4248 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.738e-13 as=1.908e-13 pd=1.79e-06 ps=1.42e-06 nrd=0.243681 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=70670 $Y=51990 $D=111
M9403 4248 4244 4245 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.738e-13 pd=1.42e-06 ps=1.79e-06 nrd=0.169811 nrs=0.243681 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=71230 $Y=51990 $D=111
M9404 4246 824 4248 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=71710 $Y=51990 $D=111
M9405 4248 824 4246 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=72190 $Y=51990 $D=111
M9406 4246 824 4248 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=1.908e-13 pd=2.76e-06 ps=1.42e-06 nrd=0.301887 nrs=0.169811 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=72670 $Y=51990 $D=111
M9407 VDD 824 4244 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.96111e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=73790 $Y=51990 $D=111
M9408 4244 824 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.89444e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=74270 $Y=51990 $D=111
M9409 VDD 824 4244 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=1.28e-06 sb=1.60574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=74750 $Y=51990 $D=111
M9410 4244 824 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.0246e-13 as=1.944e-13 pd=1.54746e-06 ps=1.44e-06 nrd=0.173577 nrs=0.166667 sa=1.76e-06 sb=1.12574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=75230 $Y=51990 $D=111
M9411 4249 4248 4244 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.7434e-13 pd=1.29e-06 ps=1.33254e-06 nrd=0.193548 nrs=0.201573 sa=2e-06 sb=7.82151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=75710 $Y=52140 $D=111
M9412 4244 4248 4249 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.81e-13 as=1.674e-13 pd=2.66e-06 ps=1.29e-06 nrd=0.324893 nrs=0.193548 sa=2e-06 sb=3.02151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=76190 $Y=52140 $D=111
M9413 4251 4247 4249 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.756e-13 pd=9.8e-07 ps=1.96e-06 nrd=0.290323 nrs=0.456816 sa=2.83226e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=77110 $Y=52310 $D=111
M9414 4249 4247 4251 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.116e-13 pd=9.8e-07 ps=9.8e-07 nrd=0.290323 nrs=0.290323 sa=7.63226e-07 sb=1.79742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=77590 $Y=52310 $D=111
M9415 4251 4247 4249 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24e-13 as=1.116e-13 pd=1.032e-06 ps=9.8e-07 nrd=0.322581 nrs=0.290323 sa=1.24323e-06 sb=1.31742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=78070 $Y=52310 $D=111
M9416 4252 4248 4251 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.86e-13 pd=1.29e-06 ps=1.548e-06 nrd=0.193548 nrs=0.215054 sa=1.24215e-06 sb=7.84946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=78550 $Y=52000 $D=111
M9417 4251 4248 4252 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.424e-13 as=1.674e-13 pd=3e-06 ps=1.29e-06 nrd=0.395884 nrs=0.193548 sa=1.58667e-06 sb=3.04946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=79030 $Y=52000 $D=111
M9418 4252 4247 4250 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=2.844e-13 pd=1.29e-06 ps=2.5e-06 nrd=0.193548 nrs=0.328824 sa=3.05806e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=80240 $Y=52210 $D=111
M9419 4250 4247 4252 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.674e-13 pd=1.29e-06 ps=1.29e-06 nrd=0.193548 nrs=0.193548 sa=7.85806e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=80720 $Y=52210 $D=111
M9420 VDD 4251 4250 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30175e-13 as=1.674e-13 pd=1.54446e-06 ps=1.29e-06 nrd=0.266129 nrs=0.193548 sa=1.26581e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=81200 $Y=52210 $D=111
M9421 4250 4251 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.296e-13 as=2.54925e-13 pd=2.7e-06 ps=1.71054e-06 nrd=0.31068 nrs=0.240291 sa=1.6835e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=81760 $Y=52110 $D=111
M9422 VDD 288 4251 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.90115e-13 as=4.128e-13 pd=1.8042e-06 ps=3.22e-06 nrd=0.174337 nrs=0.248062 sa=3.2e-07 sb=8.34419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=82700 $Y=51990 $D=111
M9423 4251 288 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.54e-13 as=2.90115e-13 pd=3.22e-06 ps=1.8042e-06 nrd=0.212728 nrs=0.174337 sa=8.8e-07 sb=2.74419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=83260 $Y=51990 $D=111
M9424 312 4249 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=84360 $Y=52000 $D=111
M9425 VDD 4249 312 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=84840 $Y=52000 $D=111
M9426 272 4252 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.56e-13 as=2.304e-13 pd=1.68e-06 ps=1.64e-06 nrd=0.15625 nrs=0.140625 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=85320 $Y=52000 $D=111
M9427 VDD 4252 272 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.56e-13 pd=3.2e-06 ps=1.68e-06 nrd=0.25 nrs=0.15625 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=85840 $Y=52000 $D=111
M9428 VDD 312 4255 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.69778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=72010 $Y=71510 $D=111
M9429 4255 312 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.21778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=72490 $Y=71510 $D=111
M9430 VDD 312 4255 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.96397e-13 as=1.944e-13 pd=1.50655e-06 ps=1.44e-06 nrd=0.168378 nrs=0.166667 sa=1.28e-06 sb=7.37778e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=72970 $Y=71510 $D=111
M9431 4253 312 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.36403e-13 pd=3.24e-06 ps=1.81345e-06 nrd=0.190769 nrs=0.139884 sa=1.496e-06 sb=2.48e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=73450 $Y=71510 $D=111
M9432 4256 4253 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=2.496e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.213992 sa=2.31111e-07 sb=1.73556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=74270 $Y=71410 $D=111
M9433 VDD 4253 4256 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=7.11111e-07 sb=1.58444e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=74750 $Y=71410 $D=111
M9434 4256 4253 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.12366e-13 as=1.944e-13 pd=1.77645e-06 ps=1.44e-06 nrd=0.18207 nrs=0.166667 sa=1.19111e-06 sb=1.43333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=75230 $Y=71410 $D=111
M9435 4257 4254 4256 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.08434e-13 pd=1.42e-06 ps=1.74355e-06 nrd=0.169811 nrs=0.185505 sa=1.25811e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=2e-15 panw7=2.08e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3.24e-14 $X=75710 $Y=71750 $D=111
M9436 4256 4254 4257 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.62264e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=76190 $Y=71750 $D=111
M9437 4257 4254 4256 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.76755e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=76670 $Y=71750 $D=111
M9438 4255 309 4257 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.91245e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=77150 $Y=71750 $D=111
M9439 4257 309 4255 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=77630 $Y=71750 $D=111
M9440 4255 309 4257 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=78110 $Y=71750 $D=111
M9441 4258 4254 4255 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=78590 $Y=71750 $D=111
M9442 4255 4254 4258 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.738e-13 as=1.908e-13 pd=1.79e-06 ps=1.42e-06 nrd=0.243681 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=79070 $Y=71750 $D=111
M9443 4258 4254 4255 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.738e-13 pd=1.42e-06 ps=1.79e-06 nrd=0.169811 nrs=0.243681 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=79630 $Y=71750 $D=111
M9444 4256 309 4258 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=80110 $Y=71750 $D=111
M9445 4258 309 4256 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=80590 $Y=71750 $D=111
M9446 4256 309 4258 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=1.908e-13 pd=2.76e-06 ps=1.42e-06 nrd=0.301887 nrs=0.169811 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=81070 $Y=71750 $D=111
M9447 VDD 309 4254 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.96111e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=82190 $Y=71730 $D=111
M9448 4254 309 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.89444e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=82670 $Y=71730 $D=111
M9449 VDD 309 4254 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=1.28e-06 sb=1.60574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=83150 $Y=71730 $D=111
M9450 4254 309 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.0246e-13 as=1.944e-13 pd=1.54746e-06 ps=1.44e-06 nrd=0.173577 nrs=0.166667 sa=1.76e-06 sb=1.12574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=83630 $Y=71730 $D=111
M9451 4259 4258 4254 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.7434e-13 pd=1.29e-06 ps=1.33254e-06 nrd=0.193548 nrs=0.201573 sa=2e-06 sb=7.82151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=84110 $Y=71730 $D=111
M9452 4254 4258 4259 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.81e-13 as=1.674e-13 pd=2.66e-06 ps=1.29e-06 nrd=0.324893 nrs=0.193548 sa=2e-06 sb=3.02151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=84590 $Y=71730 $D=111
M9453 4261 4257 4259 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.756e-13 pd=9.8e-07 ps=1.96e-06 nrd=0.290323 nrs=0.456816 sa=2.83226e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=85510 $Y=71870 $D=111
M9454 4259 4257 4261 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.116e-13 pd=9.8e-07 ps=9.8e-07 nrd=0.290323 nrs=0.290323 sa=7.63226e-07 sb=1.79742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=85990 $Y=71870 $D=111
M9455 4261 4257 4259 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24e-13 as=1.116e-13 pd=1.032e-06 ps=9.8e-07 nrd=0.322581 nrs=0.290323 sa=1.24323e-06 sb=1.31742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=86470 $Y=71870 $D=111
M9456 4262 4258 4261 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.86e-13 pd=1.29e-06 ps=1.548e-06 nrd=0.193548 nrs=0.215054 sa=1.24215e-06 sb=7.84946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=86950 $Y=71870 $D=111
M9457 4261 4258 4262 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.424e-13 as=1.674e-13 pd=3e-06 ps=1.29e-06 nrd=0.395884 nrs=0.193548 sa=1.58667e-06 sb=3.04946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=87430 $Y=71870 $D=111
M9458 4262 4257 4260 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=2.844e-13 pd=1.29e-06 ps=2.5e-06 nrd=0.193548 nrs=0.328824 sa=3.05806e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=88640 $Y=71660 $D=111
M9459 4260 4257 4262 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.674e-13 pd=1.29e-06 ps=1.29e-06 nrd=0.193548 nrs=0.193548 sa=7.85806e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=89120 $Y=71660 $D=111
M9460 VDD 4261 4260 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30175e-13 as=1.674e-13 pd=1.54446e-06 ps=1.29e-06 nrd=0.266129 nrs=0.193548 sa=1.26581e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=89600 $Y=71660 $D=111
M9461 4260 4261 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.296e-13 as=2.54925e-13 pd=2.7e-06 ps=1.71054e-06 nrd=0.31068 nrs=0.240291 sa=1.6835e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=90160 $Y=71660 $D=111
M9462 VDD 338 4261 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.90115e-13 as=4.128e-13 pd=1.8042e-06 ps=3.22e-06 nrd=0.174337 nrs=0.248062 sa=3.2e-07 sb=8.34419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=91100 $Y=71520 $D=111
M9463 4261 338 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.54e-13 as=2.90115e-13 pd=3.22e-06 ps=1.8042e-06 nrd=0.212728 nrs=0.174337 sa=8.8e-07 sb=2.74419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=91660 $Y=71520 $D=111
M9464 342 4259 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=92760 $Y=71520 $D=111
M9465 VDD 4259 342 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=93240 $Y=71520 $D=111
M9466 347 4262 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.56e-13 as=2.304e-13 pd=1.68e-06 ps=1.64e-06 nrd=0.15625 nrs=0.140625 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=93720 $Y=71520 $D=111
M9467 VDD 4262 347 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.56e-13 pd=3.2e-06 ps=1.68e-06 nrd=0.25 nrs=0.15625 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=94240 $Y=71520 $D=111
M9468 VDD 273 4265 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.69778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=72810 $Y=59410 $D=111
M9469 4265 273 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.21778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=73290 $Y=59410 $D=111
M9470 VDD 273 4265 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.96397e-13 as=1.944e-13 pd=1.50655e-06 ps=1.44e-06 nrd=0.168378 nrs=0.166667 sa=1.28e-06 sb=7.37778e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=73770 $Y=59410 $D=111
M9471 4263 273 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.36403e-13 pd=3.24e-06 ps=1.81345e-06 nrd=0.190769 nrs=0.139884 sa=1.496e-06 sb=2.48e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=74250 $Y=59190 $D=111
M9472 4266 4263 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=2.496e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.213992 sa=2.31111e-07 sb=1.73556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=75070 $Y=59510 $D=111
M9473 VDD 4263 4266 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=7.11111e-07 sb=1.58444e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=75550 $Y=59510 $D=111
M9474 4266 4263 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.12366e-13 as=1.944e-13 pd=1.77645e-06 ps=1.44e-06 nrd=0.18207 nrs=0.166667 sa=1.19111e-06 sb=1.43333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=76030 $Y=59510 $D=111
M9475 4267 4264 4266 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.08434e-13 pd=1.42e-06 ps=1.74355e-06 nrd=0.169811 nrs=0.185505 sa=1.25811e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=2e-15 panw7=2.08e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3.24e-14 $X=76510 $Y=59190 $D=111
M9476 4266 4264 4267 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.62264e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=76990 $Y=59190 $D=111
M9477 4267 4264 4266 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.76755e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=77470 $Y=59190 $D=111
M9478 4265 317 4267 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.91245e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=77950 $Y=59190 $D=111
M9479 4267 317 4265 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=78430 $Y=59190 $D=111
M9480 4265 317 4267 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=78910 $Y=59190 $D=111
M9481 4268 4264 4265 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=79390 $Y=59190 $D=111
M9482 4265 4264 4268 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.738e-13 as=1.908e-13 pd=1.79e-06 ps=1.42e-06 nrd=0.243681 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=79870 $Y=59190 $D=111
M9483 4268 4264 4265 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.738e-13 pd=1.42e-06 ps=1.79e-06 nrd=0.169811 nrs=0.243681 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=80430 $Y=59190 $D=111
M9484 4266 317 4268 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=80910 $Y=59190 $D=111
M9485 4268 317 4266 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=81390 $Y=59190 $D=111
M9486 4266 317 4268 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=1.908e-13 pd=2.76e-06 ps=1.42e-06 nrd=0.301887 nrs=0.169811 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=81870 $Y=59190 $D=111
M9487 VDD 317 4264 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.96111e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=82990 $Y=59190 $D=111
M9488 4264 317 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.89444e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=83470 $Y=59190 $D=111
M9489 VDD 317 4264 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=1.28e-06 sb=1.60574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=83950 $Y=59190 $D=111
M9490 4264 317 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.0246e-13 as=1.944e-13 pd=1.54746e-06 ps=1.44e-06 nrd=0.173577 nrs=0.166667 sa=1.76e-06 sb=1.12574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=84430 $Y=59190 $D=111
M9491 4269 4268 4264 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.7434e-13 pd=1.29e-06 ps=1.33254e-06 nrd=0.193548 nrs=0.201573 sa=2e-06 sb=7.82151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=84910 $Y=59340 $D=111
M9492 4264 4268 4269 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.81e-13 as=1.674e-13 pd=2.66e-06 ps=1.29e-06 nrd=0.324893 nrs=0.193548 sa=2e-06 sb=3.02151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=85390 $Y=59340 $D=111
M9493 4271 4267 4269 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.756e-13 pd=9.8e-07 ps=1.96e-06 nrd=0.290323 nrs=0.456816 sa=2.83226e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=86310 $Y=59510 $D=111
M9494 4269 4267 4271 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.116e-13 pd=9.8e-07 ps=9.8e-07 nrd=0.290323 nrs=0.290323 sa=7.63226e-07 sb=1.79742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=86790 $Y=59510 $D=111
M9495 4271 4267 4269 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24e-13 as=1.116e-13 pd=1.032e-06 ps=9.8e-07 nrd=0.322581 nrs=0.290323 sa=1.24323e-06 sb=1.31742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=87270 $Y=59510 $D=111
M9496 4272 4268 4271 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.86e-13 pd=1.29e-06 ps=1.548e-06 nrd=0.193548 nrs=0.215054 sa=1.24215e-06 sb=7.84946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=87750 $Y=59200 $D=111
M9497 4271 4268 4272 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.424e-13 as=1.674e-13 pd=3e-06 ps=1.29e-06 nrd=0.395884 nrs=0.193548 sa=1.58667e-06 sb=3.04946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=88230 $Y=59200 $D=111
M9498 4272 4267 4270 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=2.844e-13 pd=1.29e-06 ps=2.5e-06 nrd=0.193548 nrs=0.328824 sa=3.05806e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=89440 $Y=59410 $D=111
M9499 4270 4267 4272 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.674e-13 pd=1.29e-06 ps=1.29e-06 nrd=0.193548 nrs=0.193548 sa=7.85806e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=89920 $Y=59410 $D=111
M9500 VDD 4271 4270 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30175e-13 as=1.674e-13 pd=1.54446e-06 ps=1.29e-06 nrd=0.266129 nrs=0.193548 sa=1.26581e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=90400 $Y=59410 $D=111
M9501 4270 4271 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.296e-13 as=2.54925e-13 pd=2.7e-06 ps=1.71054e-06 nrd=0.31068 nrs=0.240291 sa=1.6835e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=90960 $Y=59310 $D=111
M9502 VDD 341 4271 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.90115e-13 as=4.128e-13 pd=1.8042e-06 ps=3.22e-06 nrd=0.174337 nrs=0.248062 sa=3.2e-07 sb=8.34419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=91900 $Y=59190 $D=111
M9503 4271 341 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.54e-13 as=2.90115e-13 pd=3.22e-06 ps=1.8042e-06 nrd=0.212728 nrs=0.174337 sa=8.8e-07 sb=2.74419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=92460 $Y=59190 $D=111
M9504 296 4269 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=93560 $Y=59200 $D=111
M9505 VDD 4269 296 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=94040 $Y=59200 $D=111
M9506 829 4272 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.56e-13 as=2.304e-13 pd=1.68e-06 ps=1.64e-06 nrd=0.15625 nrs=0.140625 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=94520 $Y=59200 $D=111
M9507 VDD 4272 829 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.56e-13 pd=3.2e-06 ps=1.68e-06 nrd=0.25 nrs=0.15625 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=95040 $Y=59200 $D=111
M9508 VDD 311 4275 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.69778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=74410 $Y=64310 $D=111
M9509 4275 311 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.21778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=74890 $Y=64310 $D=111
M9510 VDD 311 4275 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.96397e-13 as=1.944e-13 pd=1.50655e-06 ps=1.44e-06 nrd=0.168378 nrs=0.166667 sa=1.28e-06 sb=7.37778e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=75370 $Y=64310 $D=111
M9511 4273 311 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.36403e-13 pd=3.24e-06 ps=1.81345e-06 nrd=0.190769 nrs=0.139884 sa=1.496e-06 sb=2.48e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=75850 $Y=64310 $D=111
M9512 4276 4273 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=2.496e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.213992 sa=2.31111e-07 sb=1.73556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=76670 $Y=64210 $D=111
M9513 VDD 4273 4276 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=7.11111e-07 sb=1.58444e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=77150 $Y=64210 $D=111
M9514 4276 4273 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.12366e-13 as=1.944e-13 pd=1.77645e-06 ps=1.44e-06 nrd=0.18207 nrs=0.166667 sa=1.19111e-06 sb=1.43333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=77630 $Y=64210 $D=111
M9515 4277 4274 4276 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.08434e-13 pd=1.42e-06 ps=1.74355e-06 nrd=0.169811 nrs=0.185505 sa=1.25811e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=2e-15 panw7=2.08e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3.24e-14 $X=78110 $Y=64550 $D=111
M9516 4276 4274 4277 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.62264e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=78590 $Y=64550 $D=111
M9517 4277 4274 4276 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.76755e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=79070 $Y=64550 $D=111
M9518 4275 315 4277 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.91245e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=79550 $Y=64550 $D=111
M9519 4277 315 4275 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=80030 $Y=64550 $D=111
M9520 4275 315 4277 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=80510 $Y=64550 $D=111
M9521 4278 4274 4275 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=80990 $Y=64550 $D=111
M9522 4275 4274 4278 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.738e-13 as=1.908e-13 pd=1.79e-06 ps=1.42e-06 nrd=0.243681 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=81470 $Y=64550 $D=111
M9523 4278 4274 4275 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.738e-13 pd=1.42e-06 ps=1.79e-06 nrd=0.169811 nrs=0.243681 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=82030 $Y=64550 $D=111
M9524 4276 315 4278 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=82510 $Y=64550 $D=111
M9525 4278 315 4276 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=82990 $Y=64550 $D=111
M9526 4276 315 4278 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=1.908e-13 pd=2.76e-06 ps=1.42e-06 nrd=0.301887 nrs=0.169811 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=83470 $Y=64550 $D=111
M9527 VDD 315 4274 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.96111e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=84590 $Y=64530 $D=111
M9528 4274 315 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.89444e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=85070 $Y=64530 $D=111
M9529 VDD 315 4274 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=1.28e-06 sb=1.60574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=85550 $Y=64530 $D=111
M9530 4274 315 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.0246e-13 as=1.944e-13 pd=1.54746e-06 ps=1.44e-06 nrd=0.173577 nrs=0.166667 sa=1.76e-06 sb=1.12574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=86030 $Y=64530 $D=111
M9531 4279 4278 4274 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.7434e-13 pd=1.29e-06 ps=1.33254e-06 nrd=0.193548 nrs=0.201573 sa=2e-06 sb=7.82151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=86510 $Y=64530 $D=111
M9532 4274 4278 4279 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.81e-13 as=1.674e-13 pd=2.66e-06 ps=1.29e-06 nrd=0.324893 nrs=0.193548 sa=2e-06 sb=3.02151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=86990 $Y=64530 $D=111
M9533 4281 4277 4279 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.756e-13 pd=9.8e-07 ps=1.96e-06 nrd=0.290323 nrs=0.456816 sa=2.83226e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=87910 $Y=64670 $D=111
M9534 4279 4277 4281 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.116e-13 pd=9.8e-07 ps=9.8e-07 nrd=0.290323 nrs=0.290323 sa=7.63226e-07 sb=1.79742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=88390 $Y=64670 $D=111
M9535 4281 4277 4279 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24e-13 as=1.116e-13 pd=1.032e-06 ps=9.8e-07 nrd=0.322581 nrs=0.290323 sa=1.24323e-06 sb=1.31742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=88870 $Y=64670 $D=111
M9536 4282 4278 4281 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.86e-13 pd=1.29e-06 ps=1.548e-06 nrd=0.193548 nrs=0.215054 sa=1.24215e-06 sb=7.84946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=89350 $Y=64670 $D=111
M9537 4281 4278 4282 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.424e-13 as=1.674e-13 pd=3e-06 ps=1.29e-06 nrd=0.395884 nrs=0.193548 sa=1.58667e-06 sb=3.04946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=89830 $Y=64670 $D=111
M9538 4282 4277 4280 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=2.844e-13 pd=1.29e-06 ps=2.5e-06 nrd=0.193548 nrs=0.328824 sa=3.05806e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=91040 $Y=64460 $D=111
M9539 4280 4277 4282 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.674e-13 pd=1.29e-06 ps=1.29e-06 nrd=0.193548 nrs=0.193548 sa=7.85806e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=91520 $Y=64460 $D=111
M9540 VDD 4281 4280 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30175e-13 as=1.674e-13 pd=1.54446e-06 ps=1.29e-06 nrd=0.266129 nrs=0.193548 sa=1.26581e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=92000 $Y=64460 $D=111
M9541 4280 4281 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.296e-13 as=2.54925e-13 pd=2.7e-06 ps=1.71054e-06 nrd=0.31068 nrs=0.240291 sa=1.6835e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=92560 $Y=64460 $D=111
M9542 VDD 829 4281 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.90115e-13 as=4.128e-13 pd=1.8042e-06 ps=3.22e-06 nrd=0.174337 nrs=0.248062 sa=3.2e-07 sb=8.34419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=93500 $Y=64320 $D=111
M9543 4281 829 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.54e-13 as=2.90115e-13 pd=3.22e-06 ps=1.8042e-06 nrd=0.212728 nrs=0.174337 sa=8.8e-07 sb=2.74419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=94060 $Y=64320 $D=111
M9544 349 4279 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=95160 $Y=64320 $D=111
M9545 VDD 4279 349 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=95640 $Y=64320 $D=111
M9546 338 4282 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.56e-13 as=2.304e-13 pd=1.68e-06 ps=1.64e-06 nrd=0.15625 nrs=0.140625 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=96120 $Y=64320 $D=111
M9547 VDD 4282 338 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.56e-13 pd=3.2e-06 ps=1.68e-06 nrd=0.25 nrs=0.15625 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=96640 $Y=64320 $D=111
M9548 VDD 296 4285 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.69778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=77210 $Y=66610 $D=111
M9549 4285 296 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.21778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=77690 $Y=66610 $D=111
M9550 VDD 296 4285 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.96397e-13 as=1.944e-13 pd=1.50655e-06 ps=1.44e-06 nrd=0.168378 nrs=0.166667 sa=1.28e-06 sb=7.37778e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=78170 $Y=66610 $D=111
M9551 4283 296 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.36403e-13 pd=3.24e-06 ps=1.81345e-06 nrd=0.190769 nrs=0.139884 sa=1.496e-06 sb=2.48e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=78650 $Y=66390 $D=111
M9552 4286 4283 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=2.496e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.213992 sa=2.31111e-07 sb=1.73556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=79470 $Y=66710 $D=111
M9553 VDD 4283 4286 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=7.11111e-07 sb=1.58444e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=79950 $Y=66710 $D=111
M9554 4286 4283 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.12366e-13 as=1.944e-13 pd=1.77645e-06 ps=1.44e-06 nrd=0.18207 nrs=0.166667 sa=1.19111e-06 sb=1.43333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=80430 $Y=66710 $D=111
M9555 4287 4284 4286 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.08434e-13 pd=1.42e-06 ps=1.74355e-06 nrd=0.169811 nrs=0.185505 sa=1.25811e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=2e-15 panw7=2.08e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3.24e-14 $X=80910 $Y=66390 $D=111
M9556 4286 4284 4287 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.62264e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=81390 $Y=66390 $D=111
M9557 4287 4284 4286 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.76755e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=81870 $Y=66390 $D=111
M9558 4285 349 4287 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.91245e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=82350 $Y=66390 $D=111
M9559 4287 349 4285 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=82830 $Y=66390 $D=111
M9560 4285 349 4287 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=83310 $Y=66390 $D=111
M9561 4288 4284 4285 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=83790 $Y=66390 $D=111
M9562 4285 4284 4288 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.738e-13 as=1.908e-13 pd=1.79e-06 ps=1.42e-06 nrd=0.243681 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=84270 $Y=66390 $D=111
M9563 4288 4284 4285 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.738e-13 pd=1.42e-06 ps=1.79e-06 nrd=0.169811 nrs=0.243681 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=84830 $Y=66390 $D=111
M9564 4286 349 4288 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=85310 $Y=66390 $D=111
M9565 4288 349 4286 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=85790 $Y=66390 $D=111
M9566 4286 349 4288 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=1.908e-13 pd=2.76e-06 ps=1.42e-06 nrd=0.301887 nrs=0.169811 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=86270 $Y=66390 $D=111
M9567 VDD 349 4284 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.96111e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=87390 $Y=66390 $D=111
M9568 4284 349 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.89444e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=87870 $Y=66390 $D=111
M9569 VDD 349 4284 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=1.28e-06 sb=1.60574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=88350 $Y=66390 $D=111
M9570 4284 349 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.0246e-13 as=1.944e-13 pd=1.54746e-06 ps=1.44e-06 nrd=0.173577 nrs=0.166667 sa=1.76e-06 sb=1.12574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=88830 $Y=66390 $D=111
M9571 4289 4288 4284 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.7434e-13 pd=1.29e-06 ps=1.33254e-06 nrd=0.193548 nrs=0.201573 sa=2e-06 sb=7.82151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=89310 $Y=66540 $D=111
M9572 4284 4288 4289 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.81e-13 as=1.674e-13 pd=2.66e-06 ps=1.29e-06 nrd=0.324893 nrs=0.193548 sa=2e-06 sb=3.02151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=89790 $Y=66540 $D=111
M9573 4291 4287 4289 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.756e-13 pd=9.8e-07 ps=1.96e-06 nrd=0.290323 nrs=0.456816 sa=2.83226e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=90710 $Y=66710 $D=111
M9574 4289 4287 4291 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.116e-13 pd=9.8e-07 ps=9.8e-07 nrd=0.290323 nrs=0.290323 sa=7.63226e-07 sb=1.79742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=91190 $Y=66710 $D=111
M9575 4291 4287 4289 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24e-13 as=1.116e-13 pd=1.032e-06 ps=9.8e-07 nrd=0.322581 nrs=0.290323 sa=1.24323e-06 sb=1.31742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=91670 $Y=66710 $D=111
M9576 4292 4288 4291 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.86e-13 pd=1.29e-06 ps=1.548e-06 nrd=0.193548 nrs=0.215054 sa=1.24215e-06 sb=7.84946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=92150 $Y=66400 $D=111
M9577 4291 4288 4292 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.424e-13 as=1.674e-13 pd=3e-06 ps=1.29e-06 nrd=0.395884 nrs=0.193548 sa=1.58667e-06 sb=3.04946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=92630 $Y=66400 $D=111
M9578 4292 4287 4290 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=2.844e-13 pd=1.29e-06 ps=2.5e-06 nrd=0.193548 nrs=0.328824 sa=3.05806e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=93840 $Y=66610 $D=111
M9579 4290 4287 4292 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.674e-13 pd=1.29e-06 ps=1.29e-06 nrd=0.193548 nrs=0.193548 sa=7.85806e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=94320 $Y=66610 $D=111
M9580 VDD 4291 4290 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30175e-13 as=1.674e-13 pd=1.54446e-06 ps=1.29e-06 nrd=0.266129 nrs=0.193548 sa=1.26581e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=94800 $Y=66610 $D=111
M9581 4290 4291 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.296e-13 as=2.54925e-13 pd=2.7e-06 ps=1.71054e-06 nrd=0.31068 nrs=0.240291 sa=1.6835e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=95360 $Y=66510 $D=111
M9582 VDD 831 4291 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.90115e-13 as=4.128e-13 pd=1.8042e-06 ps=3.22e-06 nrd=0.174337 nrs=0.248062 sa=3.2e-07 sb=8.34419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=96300 $Y=66390 $D=111
M9583 4291 831 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.54e-13 as=2.90115e-13 pd=3.22e-06 ps=1.8042e-06 nrd=0.212728 nrs=0.174337 sa=8.8e-07 sb=2.74419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=96860 $Y=66390 $D=111
M9584 401 4289 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=97960 $Y=66400 $D=111
M9585 VDD 4289 401 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=98440 $Y=66400 $D=111
M9586 323 4292 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.56e-13 as=2.304e-13 pd=1.68e-06 ps=1.64e-06 nrd=0.15625 nrs=0.140625 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=98920 $Y=66400 $D=111
M9587 VDD 4292 323 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.56e-13 pd=3.2e-06 ps=1.68e-06 nrd=0.25 nrs=0.15625 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=99440 $Y=66400 $D=111
M9588 VDD 365 4295 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.69778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=95610 $Y=37810 $D=111
M9589 4295 365 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.21778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=96090 $Y=37810 $D=111
M9590 VDD 365 4295 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.96397e-13 as=1.944e-13 pd=1.50655e-06 ps=1.44e-06 nrd=0.168378 nrs=0.166667 sa=1.28e-06 sb=7.37778e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=96570 $Y=37810 $D=111
M9591 4293 365 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.36403e-13 pd=3.24e-06 ps=1.81345e-06 nrd=0.190769 nrs=0.139884 sa=1.496e-06 sb=2.48e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=97050 $Y=37590 $D=111
M9592 4296 4293 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=2.496e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.213992 sa=2.31111e-07 sb=1.73556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=97870 $Y=37910 $D=111
M9593 VDD 4293 4296 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=7.11111e-07 sb=1.58444e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=98350 $Y=37910 $D=111
M9594 4296 4293 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.12366e-13 as=1.944e-13 pd=1.77645e-06 ps=1.44e-06 nrd=0.18207 nrs=0.166667 sa=1.19111e-06 sb=1.43333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=98830 $Y=37910 $D=111
M9595 4297 4294 4296 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.08434e-13 pd=1.42e-06 ps=1.74355e-06 nrd=0.169811 nrs=0.185505 sa=1.25811e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=2e-15 panw7=2.08e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3.24e-14 $X=99310 $Y=37590 $D=111
M9596 4296 4294 4297 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.62264e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=99790 $Y=37590 $D=111
M9597 4297 4294 4296 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.76755e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=100270 $Y=37590 $D=111
M9598 4295 350 4297 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.91245e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=100750 $Y=37590 $D=111
M9599 4297 350 4295 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=101230 $Y=37590 $D=111
M9600 4295 350 4297 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=101710 $Y=37590 $D=111
M9601 4298 4294 4295 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=102190 $Y=37590 $D=111
M9602 4295 4294 4298 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.738e-13 as=1.908e-13 pd=1.79e-06 ps=1.42e-06 nrd=0.243681 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=102670 $Y=37590 $D=111
M9603 4298 4294 4295 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.738e-13 pd=1.42e-06 ps=1.79e-06 nrd=0.169811 nrs=0.243681 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=103230 $Y=37590 $D=111
M9604 4296 350 4298 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=103710 $Y=37590 $D=111
M9605 4298 350 4296 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=104190 $Y=37590 $D=111
M9606 4296 350 4298 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=1.908e-13 pd=2.76e-06 ps=1.42e-06 nrd=0.301887 nrs=0.169811 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=104670 $Y=37590 $D=111
M9607 VDD 350 4294 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.96111e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=105790 $Y=37590 $D=111
M9608 4294 350 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.89444e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=106270 $Y=37590 $D=111
M9609 VDD 350 4294 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=1.28e-06 sb=1.60574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=106750 $Y=37590 $D=111
M9610 4294 350 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.0246e-13 as=1.944e-13 pd=1.54746e-06 ps=1.44e-06 nrd=0.173577 nrs=0.166667 sa=1.76e-06 sb=1.12574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=107230 $Y=37590 $D=111
M9611 4299 4298 4294 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.7434e-13 pd=1.29e-06 ps=1.33254e-06 nrd=0.193548 nrs=0.201573 sa=2e-06 sb=7.82151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=107710 $Y=37740 $D=111
M9612 4294 4298 4299 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.81e-13 as=1.674e-13 pd=2.66e-06 ps=1.29e-06 nrd=0.324893 nrs=0.193548 sa=2e-06 sb=3.02151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=108190 $Y=37740 $D=111
M9613 4301 4297 4299 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.756e-13 pd=9.8e-07 ps=1.96e-06 nrd=0.290323 nrs=0.456816 sa=2.83226e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=109110 $Y=37910 $D=111
M9614 4299 4297 4301 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.116e-13 pd=9.8e-07 ps=9.8e-07 nrd=0.290323 nrs=0.290323 sa=7.63226e-07 sb=1.79742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=109590 $Y=37910 $D=111
M9615 4301 4297 4299 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24e-13 as=1.116e-13 pd=1.032e-06 ps=9.8e-07 nrd=0.322581 nrs=0.290323 sa=1.24323e-06 sb=1.31742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=110070 $Y=37910 $D=111
M9616 4302 4298 4301 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.86e-13 pd=1.29e-06 ps=1.548e-06 nrd=0.193548 nrs=0.215054 sa=1.24215e-06 sb=7.84946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=110550 $Y=37600 $D=111
M9617 4301 4298 4302 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.424e-13 as=1.674e-13 pd=3e-06 ps=1.29e-06 nrd=0.395884 nrs=0.193548 sa=1.58667e-06 sb=3.04946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=111030 $Y=37600 $D=111
M9618 4302 4297 4300 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=2.844e-13 pd=1.29e-06 ps=2.5e-06 nrd=0.193548 nrs=0.328824 sa=3.05806e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=112240 $Y=37810 $D=111
M9619 4300 4297 4302 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.674e-13 pd=1.29e-06 ps=1.29e-06 nrd=0.193548 nrs=0.193548 sa=7.85806e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=112720 $Y=37810 $D=111
M9620 VDD 4301 4300 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30175e-13 as=1.674e-13 pd=1.54446e-06 ps=1.29e-06 nrd=0.266129 nrs=0.193548 sa=1.26581e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=113200 $Y=37810 $D=111
M9621 4300 4301 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.296e-13 as=2.54925e-13 pd=2.7e-06 ps=1.71054e-06 nrd=0.31068 nrs=0.240291 sa=1.6835e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=113760 $Y=37710 $D=111
M9622 VDD 837 4301 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.90115e-13 as=4.128e-13 pd=1.8042e-06 ps=3.22e-06 nrd=0.174337 nrs=0.248062 sa=3.2e-07 sb=8.34419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=114700 $Y=37590 $D=111
M9623 4301 837 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.54e-13 as=2.90115e-13 pd=3.22e-06 ps=1.8042e-06 nrd=0.212728 nrs=0.174337 sa=8.8e-07 sb=2.74419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=115260 $Y=37590 $D=111
M9624 461 4299 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=116360 $Y=37600 $D=111
M9625 VDD 4299 461 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=116840 $Y=37600 $D=111
M9626 434 4302 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.56e-13 as=2.304e-13 pd=1.68e-06 ps=1.64e-06 nrd=0.15625 nrs=0.140625 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=117320 $Y=37600 $D=111
M9627 VDD 4302 434 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.56e-13 pd=3.2e-06 ps=1.68e-06 nrd=0.25 nrs=0.15625 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=117840 $Y=37600 $D=111
M9628 VDD 382 4305 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.69778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=100410 $Y=66610 $D=111
M9629 4305 382 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.21778e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=100890 $Y=66610 $D=111
M9630 VDD 382 4305 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.96397e-13 as=1.944e-13 pd=1.50655e-06 ps=1.44e-06 nrd=0.168378 nrs=0.166667 sa=1.28e-06 sb=7.37778e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=101370 $Y=66610 $D=111
M9631 4303 382 VDD VDD lppfet w=1.3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.224e-13 as=2.36403e-13 pd=3.24e-06 ps=1.81345e-06 nrd=0.190769 nrs=0.139884 sa=1.496e-06 sb=2.48e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=101850 $Y=66390 $D=111
M9632 4306 4303 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=2.496e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.213992 sa=2.31111e-07 sb=1.73556e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=102670 $Y=66710 $D=111
M9633 VDD 4303 4306 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=7.11111e-07 sb=1.58444e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=103150 $Y=66710 $D=111
M9634 4306 4303 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.12366e-13 as=1.944e-13 pd=1.77645e-06 ps=1.44e-06 nrd=0.18207 nrs=0.166667 sa=1.19111e-06 sb=1.43333e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.56e-14 panw10=0 $X=103630 $Y=66710 $D=111
M9635 4307 4304 4306 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.08434e-13 pd=1.42e-06 ps=1.74355e-06 nrd=0.169811 nrs=0.185505 sa=1.25811e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=2e-15 panw7=2.08e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3.24e-14 $X=104110 $Y=66390 $D=111
M9636 4306 4304 4307 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.62264e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=104590 $Y=66390 $D=111
M9637 4307 4304 4306 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.76755e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=105070 $Y=66390 $D=111
M9638 4305 434 4307 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=1.91245e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=105550 $Y=66390 $D=111
M9639 4307 434 4305 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=6e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.52e-14 $X=106030 $Y=66390 $D=111
M9640 4305 434 4307 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=106510 $Y=66390 $D=111
M9641 4308 4304 4305 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=106990 $Y=66390 $D=111
M9642 4305 4304 4308 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.738e-13 as=1.908e-13 pd=1.79e-06 ps=1.42e-06 nrd=0.243681 nrs=0.169811 sa=2e-06 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=107470 $Y=66390 $D=111
M9643 4308 4304 4305 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=2.738e-13 pd=1.42e-06 ps=1.79e-06 nrd=0.169811 nrs=0.243681 sa=2e-06 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.2e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=3e-14 $X=108030 $Y=66390 $D=111
M9644 4306 434 4308 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=108510 $Y=66390 $D=111
M9645 4308 434 4306 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.908e-13 as=1.908e-13 pd=1.42e-06 ps=1.42e-06 nrd=0.169811 nrs=0.169811 sa=2e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=108990 $Y=66390 $D=111
M9646 4306 434 4308 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.392e-13 as=1.908e-13 pd=2.76e-06 ps=1.42e-06 nrd=0.301887 nrs=0.169811 sa=2e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=109470 $Y=66390 $D=111
M9647 VDD 434 4304 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=3.456e-13 pd=1.44e-06 ps=2.8e-06 nrd=0.166667 nrs=0.296296 sa=3.2e-07 sb=1.96111e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=110590 $Y=66390 $D=111
M9648 4304 434 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=8e-07 sb=1.89444e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=111070 $Y=66390 $D=111
M9649 VDD 434 4304 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.944e-13 as=1.944e-13 pd=1.44e-06 ps=1.44e-06 nrd=0.166667 nrs=0.166667 sa=1.28e-06 sb=1.60574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=111550 $Y=66390 $D=111
M9650 4304 434 VDD VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.0246e-13 as=1.944e-13 pd=1.54746e-06 ps=1.44e-06 nrd=0.173577 nrs=0.166667 sa=1.76e-06 sb=1.12574e-06 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=6e-15 $X=112030 $Y=66390 $D=111
M9651 4309 4308 4304 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.7434e-13 pd=1.29e-06 ps=1.33254e-06 nrd=0.193548 nrs=0.201573 sa=2e-06 sb=7.82151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=112510 $Y=66540 $D=111
M9652 4304 4308 4309 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.81e-13 as=1.674e-13 pd=2.66e-06 ps=1.29e-06 nrd=0.324893 nrs=0.193548 sa=2e-06 sb=3.02151e-07 sd=0 panw1=0 panw2=0 panw3=3.6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.6e-14 panw10=0 $X=112990 $Y=66540 $D=111
M9653 4311 4307 4309 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.756e-13 pd=9.8e-07 ps=1.96e-06 nrd=0.290323 nrs=0.456816 sa=2.83226e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=113910 $Y=66710 $D=111
M9654 4309 4307 4311 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.116e-13 as=1.116e-13 pd=9.8e-07 ps=9.8e-07 nrd=0.290323 nrs=0.290323 sa=7.63226e-07 sb=1.79742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=114390 $Y=66710 $D=111
M9655 4311 4307 4309 VDD lppfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.24e-13 as=1.116e-13 pd=1.032e-06 ps=9.8e-07 nrd=0.322581 nrs=0.290323 sa=1.24323e-06 sb=1.31742e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.56e-14 panw10=0 $X=114870 $Y=66710 $D=111
M9656 4312 4308 4311 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.86e-13 pd=1.29e-06 ps=1.548e-06 nrd=0.193548 nrs=0.215054 sa=1.24215e-06 sb=7.84946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=115350 $Y=66400 $D=111
M9657 4311 4308 4312 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.424e-13 as=1.674e-13 pd=3e-06 ps=1.29e-06 nrd=0.395884 nrs=0.193548 sa=1.58667e-06 sb=3.04946e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=1.08e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=4.8e-15 $X=115830 $Y=66400 $D=111
M9658 4312 4307 4310 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=2.844e-13 pd=1.29e-06 ps=2.5e-06 nrd=0.193548 nrs=0.328824 sa=3.05806e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=117040 $Y=66610 $D=111
M9659 4310 4307 4312 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.674e-13 as=1.674e-13 pd=1.29e-06 ps=1.29e-06 nrd=0.193548 nrs=0.193548 sa=7.85806e-07 sb=1.36e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=117520 $Y=66610 $D=111
M9660 VDD 4311 4310 VDD lppfet w=9.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.30175e-13 as=1.674e-13 pd=1.54446e-06 ps=1.29e-06 nrd=0.266129 nrs=0.193548 sa=1.26581e-06 sb=8.8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.76e-14 panw10=0 $X=118000 $Y=66610 $D=111
M9661 4310 4311 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.296e-13 as=2.54925e-13 pd=2.7e-06 ps=1.71054e-06 nrd=0.31068 nrs=0.240291 sa=1.6835e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=9.6e-15 $X=118560 $Y=66510 $D=111
M9662 VDD 381 4311 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.90115e-13 as=4.128e-13 pd=1.8042e-06 ps=3.22e-06 nrd=0.174337 nrs=0.248062 sa=3.2e-07 sb=8.34419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=119500 $Y=66390 $D=111
M9663 4311 381 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.54e-13 as=2.90115e-13 pd=3.22e-06 ps=1.8042e-06 nrd=0.212728 nrs=0.174337 sa=8.8e-07 sb=2.74419e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=120060 $Y=66390 $D=111
M9664 433 4309 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.8e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=121160 $Y=66400 $D=111
M9665 VDD 4309 433 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=8e-07 sb=1.32e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=121640 $Y=66400 $D=111
M9666 392 4312 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.56e-13 as=2.304e-13 pd=1.68e-06 ps=1.64e-06 nrd=0.15625 nrs=0.140625 sa=1.28e-06 sb=8.4e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=122120 $Y=66400 $D=111
M9667 VDD 4312 392 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.56e-13 pd=3.2e-06 ps=1.68e-06 nrd=0.25 nrs=0.15625 sa=1.8e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=122640 $Y=66400 $D=111
M9668 VDD 35 4313 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.57059e-14 as=9.6e-14 pd=6.64706e-07 ps=1.24e-06 nrd=0.841176 nrs=1.06667 sa=3.2e-07 sb=1.524e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=10820 $Y=50170 $D=111
M9669 4315 13 VDD VDD lppfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37088e-13 as=1.81694e-13 pd=1.2096e-06 ps=1.59529e-06 nrd=0.264444 nrs=0.35049 sa=5.40833e-07 sb=1.64694e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=11350 $Y=50170 $D=111
M9670 28 35 4315 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.594e-13 as=1.48512e-13 pd=1.33e-06 ps=1.3104e-06 nrd=0.261999 nrs=0.244103 sa=7.83846e-07 sb=1.17256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=11830 $Y=50290 $D=111
M9671 4314 4313 28 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.106e-13 as=1.594e-13 pd=1.32e-06 ps=1.33e-06 nrd=0.346154 nrs=0.261999 sa=1.15872e-06 sb=9.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=12310 $Y=50100 $D=111
M9672 VDD 4315 4314 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=2.106e-13 pd=2.2e-06 ps=1.32e-06 nrd=0.410256 nrs=0.346154 sa=1.71026e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=12970 $Y=50100 $D=111
M9673 VDD 19 4316 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.57059e-14 as=9.6e-14 pd=6.64706e-07 ps=1.24e-06 nrd=0.841176 nrs=1.06667 sa=3.2e-07 sb=1.524e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=11220 $Y=16730 $D=111
M9674 4318 15 VDD VDD lppfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37088e-13 as=1.81694e-13 pd=1.2096e-06 ps=1.59529e-06 nrd=0.264444 nrs=0.35049 sa=5.40833e-07 sb=1.64694e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=11750 $Y=16310 $D=111
M9675 10 19 4318 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.594e-13 as=1.48512e-13 pd=1.33e-06 ps=1.3104e-06 nrd=0.261999 nrs=0.244103 sa=7.83846e-07 sb=1.17256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=12230 $Y=16130 $D=111
M9676 4317 4316 10 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.106e-13 as=1.594e-13 pd=1.32e-06 ps=1.33e-06 nrd=0.346154 nrs=0.261999 sa=1.15872e-06 sb=9.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=12710 $Y=16320 $D=111
M9677 VDD 4318 4317 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=2.106e-13 pd=2.2e-06 ps=1.32e-06 nrd=0.410256 nrs=0.346154 sa=1.71026e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=13370 $Y=16320 $D=111
M9678 VDD 802 4319 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.57059e-14 as=9.6e-14 pd=6.64706e-07 ps=1.24e-06 nrd=0.841176 nrs=1.06667 sa=3.2e-07 sb=1.524e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=18020 $Y=71770 $D=111
M9679 4321 64 VDD VDD lppfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37088e-13 as=1.81694e-13 pd=1.2096e-06 ps=1.59529e-06 nrd=0.264444 nrs=0.35049 sa=5.40833e-07 sb=1.64694e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=18550 $Y=71770 $D=111
M9680 55 802 4321 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.594e-13 as=1.48512e-13 pd=1.33e-06 ps=1.3104e-06 nrd=0.261999 nrs=0.244103 sa=7.83846e-07 sb=1.17256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=19030 $Y=71890 $D=111
M9681 4320 4319 55 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.106e-13 as=1.594e-13 pd=1.32e-06 ps=1.33e-06 nrd=0.346154 nrs=0.261999 sa=1.15872e-06 sb=9.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=19510 $Y=71700 $D=111
M9682 VDD 4321 4320 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=2.106e-13 pd=2.2e-06 ps=1.32e-06 nrd=0.410256 nrs=0.346154 sa=1.71026e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=20170 $Y=71700 $D=111
M9683 VDD 101 4322 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.57059e-14 as=9.6e-14 pd=6.64706e-07 ps=1.24e-06 nrd=0.841176 nrs=1.06667 sa=3.2e-07 sb=1.524e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=26020 $Y=28570 $D=111
M9684 4324 78 VDD VDD lppfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37088e-13 as=1.81694e-13 pd=1.2096e-06 ps=1.59529e-06 nrd=0.264444 nrs=0.35049 sa=5.40833e-07 sb=1.64694e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=26550 $Y=28570 $D=111
M9685 83 101 4324 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.594e-13 as=1.48512e-13 pd=1.33e-06 ps=1.3104e-06 nrd=0.261999 nrs=0.244103 sa=7.83846e-07 sb=1.17256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=27030 $Y=28690 $D=111
M9686 4323 4322 83 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.106e-13 as=1.594e-13 pd=1.32e-06 ps=1.33e-06 nrd=0.346154 nrs=0.261999 sa=1.15872e-06 sb=9.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=27510 $Y=28500 $D=111
M9687 VDD 4324 4323 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=2.106e-13 pd=2.2e-06 ps=1.32e-06 nrd=0.410256 nrs=0.346154 sa=1.71026e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=28170 $Y=28500 $D=111
M9688 VDD 163 4325 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.57059e-14 as=9.6e-14 pd=6.64706e-07 ps=1.24e-06 nrd=0.841176 nrs=1.06667 sa=3.2e-07 sb=1.524e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=46820 $Y=31130 $D=111
M9689 4327 176 VDD VDD lppfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37088e-13 as=1.81694e-13 pd=1.2096e-06 ps=1.59529e-06 nrd=0.264444 nrs=0.35049 sa=5.40833e-07 sb=1.64694e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=47350 $Y=30710 $D=111
M9690 164 163 4327 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.594e-13 as=1.48512e-13 pd=1.33e-06 ps=1.3104e-06 nrd=0.261999 nrs=0.244103 sa=7.83846e-07 sb=1.17256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=47830 $Y=30530 $D=111
M9691 4326 4325 164 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.106e-13 as=1.594e-13 pd=1.32e-06 ps=1.33e-06 nrd=0.346154 nrs=0.261999 sa=1.15872e-06 sb=9.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=48310 $Y=30720 $D=111
M9692 VDD 4327 4326 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=2.106e-13 pd=2.2e-06 ps=1.32e-06 nrd=0.410256 nrs=0.346154 sa=1.71026e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=48970 $Y=30720 $D=111
M9693 VDD 114 4328 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.57059e-14 as=9.6e-14 pd=6.64706e-07 ps=1.24e-06 nrd=0.841176 nrs=1.06667 sa=3.2e-07 sb=1.524e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=48820 $Y=50170 $D=111
M9694 4330 183 VDD VDD lppfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37088e-13 as=1.81694e-13 pd=1.2096e-06 ps=1.59529e-06 nrd=0.264444 nrs=0.35049 sa=5.40833e-07 sb=1.64694e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=49350 $Y=50170 $D=111
M9695 185 114 4330 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.594e-13 as=1.48512e-13 pd=1.33e-06 ps=1.3104e-06 nrd=0.261999 nrs=0.244103 sa=7.83846e-07 sb=1.17256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=49830 $Y=50290 $D=111
M9696 4329 4328 185 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.106e-13 as=1.594e-13 pd=1.32e-06 ps=1.33e-06 nrd=0.346154 nrs=0.261999 sa=1.15872e-06 sb=9.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=50310 $Y=50100 $D=111
M9697 VDD 4330 4329 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=2.106e-13 pd=2.2e-06 ps=1.32e-06 nrd=0.410256 nrs=0.346154 sa=1.71026e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=50970 $Y=50100 $D=111
M9698 VDD 114 4331 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.57059e-14 as=9.6e-14 pd=6.64706e-07 ps=1.24e-06 nrd=0.841176 nrs=1.06667 sa=3.2e-07 sb=1.524e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=50020 $Y=57370 $D=111
M9699 4333 186 VDD VDD lppfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37088e-13 as=1.81694e-13 pd=1.2096e-06 ps=1.59529e-06 nrd=0.264444 nrs=0.35049 sa=5.40833e-07 sb=1.64694e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=50550 $Y=57370 $D=111
M9700 200 114 4333 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.594e-13 as=1.48512e-13 pd=1.33e-06 ps=1.3104e-06 nrd=0.261999 nrs=0.244103 sa=7.83846e-07 sb=1.17256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=51030 $Y=57490 $D=111
M9701 4332 4331 200 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.106e-13 as=1.594e-13 pd=1.32e-06 ps=1.33e-06 nrd=0.346154 nrs=0.261999 sa=1.15872e-06 sb=9.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=51510 $Y=57300 $D=111
M9702 VDD 4333 4332 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=2.106e-13 pd=2.2e-06 ps=1.32e-06 nrd=0.410256 nrs=0.346154 sa=1.71026e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=52170 $Y=57300 $D=111
M9703 VDD 816 4334 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.57059e-14 as=9.6e-14 pd=6.64706e-07 ps=1.24e-06 nrd=0.841176 nrs=1.06667 sa=3.2e-07 sb=1.524e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=58020 $Y=21370 $D=111
M9704 4336 235 VDD VDD lppfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37088e-13 as=1.81694e-13 pd=1.2096e-06 ps=1.59529e-06 nrd=0.264444 nrs=0.35049 sa=5.40833e-07 sb=1.64694e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=58550 $Y=21370 $D=111
M9705 817 816 4336 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.594e-13 as=1.48512e-13 pd=1.33e-06 ps=1.3104e-06 nrd=0.261999 nrs=0.244103 sa=7.83846e-07 sb=1.17256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=59030 $Y=21490 $D=111
M9706 4335 4334 817 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.106e-13 as=1.594e-13 pd=1.32e-06 ps=1.33e-06 nrd=0.346154 nrs=0.261999 sa=1.15872e-06 sb=9.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=59510 $Y=21300 $D=111
M9707 VDD 4336 4335 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=2.106e-13 pd=2.2e-06 ps=1.32e-06 nrd=0.410256 nrs=0.346154 sa=1.71026e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=60170 $Y=21300 $D=111
M9708 VDD 228 4337 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.57059e-14 as=9.6e-14 pd=6.64706e-07 ps=1.24e-06 nrd=0.841176 nrs=1.06667 sa=3.2e-07 sb=1.524e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=68020 $Y=50170 $D=111
M9709 4339 283 VDD VDD lppfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37088e-13 as=1.81694e-13 pd=1.2096e-06 ps=1.59529e-06 nrd=0.264444 nrs=0.35049 sa=5.40833e-07 sb=1.64694e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=68550 $Y=50170 $D=111
M9710 255 228 4339 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.594e-13 as=1.48512e-13 pd=1.33e-06 ps=1.3104e-06 nrd=0.261999 nrs=0.244103 sa=7.83846e-07 sb=1.17256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=69030 $Y=50290 $D=111
M9711 4338 4337 255 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.106e-13 as=1.594e-13 pd=1.32e-06 ps=1.33e-06 nrd=0.346154 nrs=0.261999 sa=1.15872e-06 sb=9.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=69510 $Y=50100 $D=111
M9712 VDD 4339 4338 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=2.106e-13 pd=2.2e-06 ps=1.32e-06 nrd=0.410256 nrs=0.346154 sa=1.71026e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=70170 $Y=50100 $D=111
M9713 VDD 411 4340 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.57059e-14 as=9.6e-14 pd=6.64706e-07 ps=1.24e-06 nrd=0.841176 nrs=1.06667 sa=3.2e-07 sb=1.524e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=7.2e-15 panw9=0 panw10=0 $X=100020 $Y=64570 $D=111
M9714 4342 372 VDD VDD lppfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.37088e-13 as=1.81694e-13 pd=1.2096e-06 ps=1.59529e-06 nrd=0.264444 nrs=0.35049 sa=5.40833e-07 sb=1.64694e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=4.8e-15 panw7=2.4e-14 panw8=2.4e-14 panw9=3.36e-14 panw10=0 $X=100550 $Y=64570 $D=111
M9715 370 411 4342 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.594e-13 as=1.48512e-13 pd=1.33e-06 ps=1.3104e-06 nrd=0.261999 nrs=0.244103 sa=7.83846e-07 sb=1.17256e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.44e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=7.2e-15 $X=101030 $Y=64690 $D=111
M9716 4341 4340 370 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.106e-13 as=1.594e-13 pd=1.32e-06 ps=1.33e-06 nrd=0.346154 nrs=0.261999 sa=1.15872e-06 sb=9.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=101510 $Y=64500 $D=111
M9717 VDD 4342 4341 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.496e-13 as=2.106e-13 pd=2.2e-06 ps=1.32e-06 nrd=0.410256 nrs=0.346154 sa=1.71026e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=1.2e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.24e-14 panw10=0 $X=102170 $Y=64500 $D=111
M9718 4343 73 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.854e-13 as=3.296e-13 pd=1.39e-06 ps=2.7e-06 nrd=0.174757 nrs=0.31068 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=23210 $Y=57120 $D=111
M9719 VDD 73 4343 VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8755e-13 as=1.854e-13 pd=1.45991e-06 ps=1.39e-06 nrd=0.176783 nrs=0.174757 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=23690 $Y=57120 $D=111
M9720 82 4343 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.3125e-13 pd=1.63e-06 ps=1.80009e-06 nrd=0.141732 nrs=0.143376 sa=1.07591e-06 sb=1.84e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=24170 $Y=57120 $D=111
M9721 VDD 4343 82 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.86913e-13 as=2.286e-13 pd=1.78873e-06 ps=1.63e-06 nrd=0.177886 nrs=0.141732 sa=1.55591e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=24650 $Y=57120 $D=111
M9722 82 4343 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.91431e-13 pd=1.65e-06 ps=1.8169e-06 nrd=0.139535 nrs=0.175128 sa=1.83318e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=25210 $Y=57120 $D=111
M9723 VDD 4343 82 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=1.92992e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=25690 $Y=57120 $D=111
M9724 4344 98 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.854e-13 as=3.296e-13 pd=1.39e-06 ps=2.7e-06 nrd=0.174757 nrs=0.31068 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=23610 $Y=42720 $D=111
M9725 VDD 98 4344 VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8755e-13 as=1.854e-13 pd=1.45991e-06 ps=1.39e-06 nrd=0.176783 nrs=0.174757 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=24090 $Y=42720 $D=111
M9726 84 4344 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.3125e-13 pd=1.63e-06 ps=1.80009e-06 nrd=0.141732 nrs=0.143376 sa=1.07591e-06 sb=1.84e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=24570 $Y=42720 $D=111
M9727 VDD 4344 84 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.86913e-13 as=2.286e-13 pd=1.78873e-06 ps=1.63e-06 nrd=0.177886 nrs=0.141732 sa=1.55591e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=25050 $Y=42720 $D=111
M9728 84 4344 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.91431e-13 pd=1.65e-06 ps=1.8169e-06 nrd=0.139535 nrs=0.175128 sa=1.83318e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=25610 $Y=42720 $D=111
M9729 VDD 4344 84 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=1.92992e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=26090 $Y=42720 $D=111
M9730 4345 114 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.854e-13 as=3.296e-13 pd=1.39e-06 ps=2.7e-06 nrd=0.174757 nrs=0.31068 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=31610 $Y=28320 $D=111
M9731 VDD 114 4345 VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8755e-13 as=1.854e-13 pd=1.45991e-06 ps=1.39e-06 nrd=0.176783 nrs=0.174757 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=32090 $Y=28320 $D=111
M9732 113 4345 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.3125e-13 pd=1.63e-06 ps=1.80009e-06 nrd=0.141732 nrs=0.143376 sa=1.07591e-06 sb=1.84e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=32570 $Y=28320 $D=111
M9733 VDD 4345 113 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.86913e-13 as=2.286e-13 pd=1.78873e-06 ps=1.63e-06 nrd=0.177886 nrs=0.141732 sa=1.55591e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=33050 $Y=28320 $D=111
M9734 113 4345 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.91431e-13 pd=1.65e-06 ps=1.8169e-06 nrd=0.139535 nrs=0.175128 sa=1.83318e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=33610 $Y=28320 $D=111
M9735 VDD 4345 113 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=1.92992e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=34090 $Y=28320 $D=111
M9736 4346 111 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.854e-13 as=3.296e-13 pd=1.39e-06 ps=2.7e-06 nrd=0.174757 nrs=0.31068 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=33210 $Y=73850 $D=111
M9737 VDD 111 4346 VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8755e-13 as=1.854e-13 pd=1.45991e-06 ps=1.39e-06 nrd=0.176783 nrs=0.174757 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=33690 $Y=73850 $D=111
M9738 89 4346 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.3125e-13 pd=1.63e-06 ps=1.80009e-06 nrd=0.141732 nrs=0.143376 sa=1.07591e-06 sb=1.84e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=34170 $Y=73610 $D=111
M9739 VDD 4346 89 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.86913e-13 as=2.286e-13 pd=1.78873e-06 ps=1.63e-06 nrd=0.177886 nrs=0.141732 sa=1.55591e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=34650 $Y=73610 $D=111
M9740 89 4346 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.91431e-13 pd=1.65e-06 ps=1.8169e-06 nrd=0.139535 nrs=0.175128 sa=1.83318e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=35210 $Y=73590 $D=111
M9741 VDD 4346 89 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=1.92992e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=35690 $Y=73590 $D=111
M9742 4347 136 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.854e-13 as=3.296e-13 pd=1.39e-06 ps=2.7e-06 nrd=0.174757 nrs=0.31068 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=37210 $Y=45050 $D=111
M9743 VDD 136 4347 VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8755e-13 as=1.854e-13 pd=1.45991e-06 ps=1.39e-06 nrd=0.176783 nrs=0.174757 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=37690 $Y=45050 $D=111
M9744 176 4347 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.3125e-13 pd=1.63e-06 ps=1.80009e-06 nrd=0.141732 nrs=0.143376 sa=1.07591e-06 sb=1.84e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=38170 $Y=44810 $D=111
M9745 VDD 4347 176 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.86913e-13 as=2.286e-13 pd=1.78873e-06 ps=1.63e-06 nrd=0.177886 nrs=0.141732 sa=1.55591e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=38650 $Y=44810 $D=111
M9746 176 4347 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.91431e-13 pd=1.65e-06 ps=1.8169e-06 nrd=0.139535 nrs=0.175128 sa=1.83318e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=39210 $Y=44790 $D=111
M9747 VDD 4347 176 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=1.92992e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=39690 $Y=44790 $D=111
M9748 4348 129 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.854e-13 as=3.296e-13 pd=1.39e-06 ps=2.7e-06 nrd=0.174757 nrs=0.31068 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=49610 $Y=42720 $D=111
M9749 VDD 129 4348 VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8755e-13 as=1.854e-13 pd=1.45991e-06 ps=1.39e-06 nrd=0.176783 nrs=0.174757 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=50090 $Y=42720 $D=111
M9750 228 4348 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.3125e-13 pd=1.63e-06 ps=1.80009e-06 nrd=0.141732 nrs=0.143376 sa=1.07591e-06 sb=1.84e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=50570 $Y=42720 $D=111
M9751 VDD 4348 228 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.86913e-13 as=2.286e-13 pd=1.78873e-06 ps=1.63e-06 nrd=0.177886 nrs=0.141732 sa=1.55591e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=51050 $Y=42720 $D=111
M9752 228 4348 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.91431e-13 pd=1.65e-06 ps=1.8169e-06 nrd=0.139535 nrs=0.175128 sa=1.83318e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=51610 $Y=42720 $D=111
M9753 VDD 4348 228 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=1.92992e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=52090 $Y=42720 $D=111
M9754 4349 283 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.854e-13 as=3.296e-13 pd=1.39e-06 ps=2.7e-06 nrd=0.174757 nrs=0.31068 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=75610 $Y=45050 $D=111
M9755 VDD 283 4349 VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8755e-13 as=1.854e-13 pd=1.45991e-06 ps=1.39e-06 nrd=0.176783 nrs=0.174757 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=76090 $Y=45050 $D=111
M9756 354 4349 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.3125e-13 pd=1.63e-06 ps=1.80009e-06 nrd=0.141732 nrs=0.143376 sa=1.07591e-06 sb=1.84e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=76570 $Y=44810 $D=111
M9757 VDD 4349 354 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.86913e-13 as=2.286e-13 pd=1.78873e-06 ps=1.63e-06 nrd=0.177886 nrs=0.141732 sa=1.55591e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=77050 $Y=44810 $D=111
M9758 354 4349 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.91431e-13 pd=1.65e-06 ps=1.8169e-06 nrd=0.139535 nrs=0.175128 sa=1.83318e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=77610 $Y=44790 $D=111
M9759 VDD 4349 354 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=1.92992e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=78090 $Y=44790 $D=111
M9760 4350 354 VDD VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.854e-13 as=3.296e-13 pd=1.39e-06 ps=2.7e-06 nrd=0.174757 nrs=0.31068 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=98810 $Y=49920 $D=111
M9761 VDD 354 4350 VDD lppfet w=1.03e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.8755e-13 as=1.854e-13 pd=1.45991e-06 ps=1.39e-06 nrd=0.176783 nrs=0.174757 sa=8e-07 sb=2e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.08e-14 panw10=0 $X=99290 $Y=49920 $D=111
M9762 395 4350 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.3125e-13 pd=1.63e-06 ps=1.80009e-06 nrd=0.141732 nrs=0.143376 sa=1.07591e-06 sb=1.84e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=99770 $Y=49920 $D=111
M9763 VDD 4350 395 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.86913e-13 as=2.286e-13 pd=1.78873e-06 ps=1.63e-06 nrd=0.177886 nrs=0.141732 sa=1.55591e-06 sb=1.36e-06 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=100250 $Y=49920 $D=111
M9764 395 4350 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.91431e-13 pd=1.65e-06 ps=1.8169e-06 nrd=0.139535 nrs=0.175128 sa=1.83318e-06 sb=8e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=100810 $Y=49920 $D=111
M9765 VDD 4350 395 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.128e-13 as=2.322e-13 pd=3.22e-06 ps=1.65e-06 nrd=0.248062 nrs=0.139535 sa=1.92992e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=101290 $Y=49920 $D=111
M9766 4351 86 VDD VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=2.464e-13 pd=1.13e-06 ps=2.18e-06 nrd=0.233766 nrs=0.415584 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=28660 $Y=57110 $D=111
M9767 VDD 86 4351 VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.70453e-13 as=1.386e-13 pd=1.32282e-06 ps=1.13e-06 nrd=0.28749 nrs=0.233766 sa=8e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=29140 $Y=57110 $D=111
M9768 114 4351 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.85564e-13 pd=1.65e-06 ps=2.21615e-06 nrd=0.139535 nrs=0.171603 sa=8.89922e-07 sb=1.34791e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=29620 $Y=57110 $D=111
M9769 VDD 4351 114 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93372e-13 as=2.322e-13 pd=1.83244e-06 ps=1.65e-06 nrd=0.176295 nrs=0.139535 sa=1.36992e-06 sb=8.67907e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=30100 $Y=57110 $D=111
M9770 114 4351 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.032e-13 as=2.8655e-13 pd=3.16e-06 ps=1.78982e-06 nrd=0.253968 nrs=0.180492 sa=1.74698e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=30660 $Y=57110 $D=111
M9771 4352 89 VDD VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=2.464e-13 pd=1.13e-06 ps=2.18e-06 nrd=0.233766 nrs=0.415584 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=30260 $Y=74120 $D=111
M9772 VDD 89 4352 VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.70453e-13 as=1.386e-13 pd=1.32282e-06 ps=1.13e-06 nrd=0.28749 nrs=0.233766 sa=8e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=30740 $Y=74120 $D=111
M9773 162 4352 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.85564e-13 pd=1.65e-06 ps=2.21615e-06 nrd=0.139535 nrs=0.171603 sa=8.89922e-07 sb=1.34791e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=31220 $Y=73600 $D=111
M9774 VDD 4352 162 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93372e-13 as=2.322e-13 pd=1.83244e-06 ps=1.65e-06 nrd=0.176295 nrs=0.139535 sa=1.36992e-06 sb=8.67907e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=31700 $Y=73600 $D=111
M9775 162 4352 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.032e-13 as=2.8655e-13 pd=3.16e-06 ps=1.78982e-06 nrd=0.253968 nrs=0.180492 sa=1.74698e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=32260 $Y=73630 $D=111
M9776 4353 114 VDD VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=2.464e-13 pd=1.13e-06 ps=2.18e-06 nrd=0.233766 nrs=0.415584 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=37060 $Y=49910 $D=111
M9777 VDD 114 4353 VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.70453e-13 as=1.386e-13 pd=1.32282e-06 ps=1.13e-06 nrd=0.28749 nrs=0.233766 sa=8e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=37540 $Y=49910 $D=111
M9778 163 4353 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.85564e-13 pd=1.65e-06 ps=2.21615e-06 nrd=0.139535 nrs=0.171603 sa=8.89922e-07 sb=1.34791e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=38020 $Y=49910 $D=111
M9779 VDD 4353 163 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93372e-13 as=2.322e-13 pd=1.83244e-06 ps=1.65e-06 nrd=0.176295 nrs=0.139535 sa=1.36992e-06 sb=8.67907e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=38500 $Y=49910 $D=111
M9780 163 4353 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.032e-13 as=2.8655e-13 pd=3.16e-06 ps=1.78982e-06 nrd=0.253968 nrs=0.180492 sa=1.74698e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=39060 $Y=49910 $D=111
M9781 4354 894 VDD VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=2.464e-13 pd=1.13e-06 ps=2.18e-06 nrd=0.233766 nrs=0.415584 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=48260 $Y=64310 $D=111
M9782 VDD 894 4354 VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.70453e-13 as=1.386e-13 pd=1.32282e-06 ps=1.13e-06 nrd=0.28749 nrs=0.233766 sa=8e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=48740 $Y=64310 $D=111
M9783 248 4354 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.85564e-13 pd=1.65e-06 ps=2.21615e-06 nrd=0.139535 nrs=0.171603 sa=8.89922e-07 sb=1.34791e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=49220 $Y=64310 $D=111
M9784 VDD 4354 248 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93372e-13 as=2.322e-13 pd=1.83244e-06 ps=1.65e-06 nrd=0.176295 nrs=0.139535 sa=1.36992e-06 sb=8.67907e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=49700 $Y=64310 $D=111
M9785 248 4354 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.032e-13 as=2.8655e-13 pd=3.16e-06 ps=1.78982e-06 nrd=0.253968 nrs=0.180492 sa=1.74698e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=50260 $Y=64310 $D=111
M9786 4355 182 VDD VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=2.464e-13 pd=1.13e-06 ps=2.18e-06 nrd=0.233766 nrs=0.415584 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=49460 $Y=23720 $D=111
M9787 VDD 182 4355 VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.70453e-13 as=1.386e-13 pd=1.32282e-06 ps=1.13e-06 nrd=0.28749 nrs=0.233766 sa=8e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=49940 $Y=23720 $D=111
M9788 198 4355 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.85564e-13 pd=1.65e-06 ps=2.21615e-06 nrd=0.139535 nrs=0.171603 sa=8.89922e-07 sb=1.34791e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=50420 $Y=23200 $D=111
M9789 VDD 4355 198 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93372e-13 as=2.322e-13 pd=1.83244e-06 ps=1.65e-06 nrd=0.176295 nrs=0.139535 sa=1.36992e-06 sb=8.67907e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=50900 $Y=23200 $D=111
M9790 198 4355 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.032e-13 as=2.8655e-13 pd=3.16e-06 ps=1.78982e-06 nrd=0.253968 nrs=0.180492 sa=1.74698e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=51460 $Y=23230 $D=111
M9791 4356 213 VDD VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=2.464e-13 pd=1.13e-06 ps=2.18e-06 nrd=0.233766 nrs=0.415584 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=71460 $Y=49910 $D=111
M9792 VDD 213 4356 VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.70453e-13 as=1.386e-13 pd=1.32282e-06 ps=1.13e-06 nrd=0.28749 nrs=0.233766 sa=8e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=71940 $Y=49910 $D=111
M9793 325 4356 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.85564e-13 pd=1.65e-06 ps=2.21615e-06 nrd=0.139535 nrs=0.171603 sa=8.89922e-07 sb=1.34791e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=72420 $Y=49910 $D=111
M9794 VDD 4356 325 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93372e-13 as=2.322e-13 pd=1.83244e-06 ps=1.65e-06 nrd=0.176295 nrs=0.139535 sa=1.36992e-06 sb=8.67907e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=72900 $Y=49910 $D=111
M9795 325 4356 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.032e-13 as=2.8655e-13 pd=3.16e-06 ps=1.78982e-06 nrd=0.253968 nrs=0.180492 sa=1.74698e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=73460 $Y=49910 $D=111
M9796 4357 320 VDD VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=2.464e-13 pd=1.13e-06 ps=2.18e-06 nrd=0.233766 nrs=0.415584 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=81060 $Y=49910 $D=111
M9797 VDD 320 4357 VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.70453e-13 as=1.386e-13 pd=1.32282e-06 ps=1.13e-06 nrd=0.28749 nrs=0.233766 sa=8e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=81540 $Y=49910 $D=111
M9798 311 4357 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.85564e-13 pd=1.65e-06 ps=2.21615e-06 nrd=0.139535 nrs=0.171603 sa=8.89922e-07 sb=1.34791e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=82020 $Y=49910 $D=111
M9799 VDD 4357 311 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93372e-13 as=2.322e-13 pd=1.83244e-06 ps=1.65e-06 nrd=0.176295 nrs=0.139535 sa=1.36992e-06 sb=8.67907e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=82500 $Y=49910 $D=111
M9800 311 4357 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.032e-13 as=2.8655e-13 pd=3.16e-06 ps=1.78982e-06 nrd=0.253968 nrs=0.180492 sa=1.74698e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=83060 $Y=49910 $D=111
M9801 4358 346 VDD VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=2.464e-13 pd=1.13e-06 ps=2.18e-06 nrd=0.233766 nrs=0.415584 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=83060 $Y=38120 $D=111
M9802 VDD 346 4358 VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.70453e-13 as=1.386e-13 pd=1.32282e-06 ps=1.13e-06 nrd=0.28749 nrs=0.233766 sa=8e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=83540 $Y=38120 $D=111
M9803 350 4358 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.85564e-13 pd=1.65e-06 ps=2.21615e-06 nrd=0.139535 nrs=0.171603 sa=8.89922e-07 sb=1.34791e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=84020 $Y=37600 $D=111
M9804 VDD 4358 350 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93372e-13 as=2.322e-13 pd=1.83244e-06 ps=1.65e-06 nrd=0.176295 nrs=0.139535 sa=1.36992e-06 sb=8.67907e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=84500 $Y=37600 $D=111
M9805 350 4358 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.032e-13 as=2.8655e-13 pd=3.16e-06 ps=1.78982e-06 nrd=0.253968 nrs=0.180492 sa=1.74698e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=85060 $Y=37630 $D=111
M9806 4359 325 VDD VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=2.464e-13 pd=1.13e-06 ps=2.18e-06 nrd=0.233766 nrs=0.415584 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=89860 $Y=45320 $D=111
M9807 VDD 325 4359 VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.70453e-13 as=1.386e-13 pd=1.32282e-06 ps=1.13e-06 nrd=0.28749 nrs=0.233766 sa=8e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=90340 $Y=45320 $D=111
M9808 400 4359 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.85564e-13 pd=1.65e-06 ps=2.21615e-06 nrd=0.139535 nrs=0.171603 sa=8.89922e-07 sb=1.34791e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=90820 $Y=44800 $D=111
M9809 VDD 4359 400 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93372e-13 as=2.322e-13 pd=1.83244e-06 ps=1.65e-06 nrd=0.176295 nrs=0.139535 sa=1.36992e-06 sb=8.67907e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=91300 $Y=44800 $D=111
M9810 400 4359 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.032e-13 as=2.8655e-13 pd=3.16e-06 ps=1.78982e-06 nrd=0.253968 nrs=0.180492 sa=1.74698e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=91860 $Y=44830 $D=111
M9811 4360 246 VDD VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.386e-13 as=2.464e-13 pd=1.13e-06 ps=2.18e-06 nrd=0.233766 nrs=0.415584 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=93060 $Y=45320 $D=111
M9812 VDD 246 4360 VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.70453e-13 as=1.386e-13 pd=1.32282e-06 ps=1.13e-06 nrd=0.28749 nrs=0.233766 sa=8e-07 sb=1.84e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=93540 $Y=45320 $D=111
M9813 410 4360 VDD VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.322e-13 as=2.85564e-13 pd=1.65e-06 ps=2.21615e-06 nrd=0.139535 nrs=0.171603 sa=8.89922e-07 sb=1.34791e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=94020 $Y=44800 $D=111
M9814 VDD 4360 410 VDD lppfet w=1.29e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.93372e-13 as=2.322e-13 pd=1.83244e-06 ps=1.65e-06 nrd=0.176295 nrs=0.139535 sa=1.36992e-06 sb=8.67907e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.28e-14 $X=94500 $Y=44800 $D=111
M9815 410 4360 VDD VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.032e-13 as=2.8655e-13 pd=3.16e-06 ps=1.78982e-06 nrd=0.253968 nrs=0.180492 sa=1.74698e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.92e-14 $X=95060 $Y=44830 $D=111
M9816 291 284 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=76010 $Y=35510 $D=111
M9817 VDD 284 291 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8791e-13 as=2.304e-13 pd=1.7938e-06 ps=1.64e-06 nrd=0.175726 nrs=0.140625 sa=8e-07 sb=8.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=76490 $Y=35510 $D=111
M9818 291 284 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.224e-13 as=2.8791e-13 pd=3.22e-06 ps=1.7938e-06 nrd=0.257812 nrs=0.175726 sa=1.36e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=77050 $Y=35510 $D=111
M9819 304 284 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=78010 $Y=35510 $D=111
M9820 VDD 284 304 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8791e-13 as=2.304e-13 pd=1.7938e-06 ps=1.64e-06 nrd=0.175726 nrs=0.140625 sa=8e-07 sb=8.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=78490 $Y=35510 $D=111
M9821 304 284 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.224e-13 as=2.8791e-13 pd=3.22e-06 ps=1.7938e-06 nrd=0.257812 nrs=0.175726 sa=1.36e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=79050 $Y=35510 $D=111
M9822 316 302 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.37e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=84010 $Y=13910 $D=111
M9823 VDD 302 316 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8791e-13 as=2.304e-13 pd=1.7938e-06 ps=1.64e-06 nrd=0.175726 nrs=0.140625 sa=8e-07 sb=8.9e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=84490 $Y=13910 $D=111
M9824 316 302 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.224e-13 as=2.8791e-13 pd=3.22e-06 ps=1.7938e-06 nrd=0.257812 nrs=0.175726 sa=1.36e-06 sb=3.3e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=85050 $Y=13910 $D=111
M9825 265 242 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.304e-13 pd=1.92e-06 ps=2e-06 nrd=0.5 nrs=0.5625 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=68570 $Y=45450 $D=111
M9826 297 313 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=2.304e-13 pd=1.92e-06 ps=2e-06 nrd=0.5 nrs=0.5625 sa=3.6e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=78570 $Y=42710 $D=111
M9827 4370 798 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=12860 $Y=14640 $D=111
M9828 4362 4364 4370 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=13180 $Y=14640 $D=111
M9829 VDD 76 4362 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=13660 $Y=14640 $D=111
M9830 VDD clk 4361 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=14180 $Y=13910 $D=111
M9831 4364 4361 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=14690 $Y=13910 $D=111
M9832 4372 4361 4362 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=15250 $Y=14410 $D=111
M9833 VDD 4363 4372 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=15570 $Y=14410 $D=111
M9834 4363 4362 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=16110 $Y=14410 $D=111
M9835 4365 4361 4363 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.83893e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.16e-14 panw9=1.2e-14 panw10=0 $X=16940 $Y=14660 $D=111
M9836 4375 4364 4365 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=1.41857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.16e-14 panw9=1.2e-14 panw10=0 $X=17670 $Y=14660 $D=111
M9837 VDD 4368 4375 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30238e-13 as=2.94e-14 pd=8.27387e-07 ps=4.9e-07 nrd=1.6612 nrs=0.375 sa=1.72321e-06 sb=1.08857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=18000 $Y=14660 $D=111
M9838 4368 76 VDD VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.84e-14 as=1.76751e-13 pd=7.4e-07 ps=1.12288e-06 nrd=0.473684 nrs=1.22404 sa=1.18763e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=2.64e-14 panw10=0 $X=18730 $Y=14450 $D=111
M9839 VDD 4365 4368 VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50686e-13 as=6.84e-14 pd=1.39215e-06 ps=7.4e-07 nrd=1.04353 nrs=0.473684 sa=1.45289e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=2.64e-14 panw10=0 $X=19210 $Y=14450 $D=111
M9840 4366 4368 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.18963e-13 pd=1.24e-06 ps=1.09907e-06 nrd=1.06667 nrs=1.32181 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=19650 $Y=14050 $D=111
M9841 VDD 4366 4367 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=20590 $Y=13930 $D=111
M9842 62 4368 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=21070 $Y=13930 $D=111
M9843 4387 24 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=16060 $Y=59480 $D=111
M9844 4379 4381 4387 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=16380 $Y=59480 $D=111
M9845 VDD 32 4379 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=16860 $Y=59480 $D=111
M9846 VDD clk 4378 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=17380 $Y=60070 $D=111
M9847 4381 4378 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=17890 $Y=60210 $D=111
M9848 4389 4378 4379 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=18450 $Y=59710 $D=111
M9849 VDD 4380 4389 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=18770 $Y=59710 $D=111
M9850 4380 4379 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=19310 $Y=59710 $D=111
M9851 4382 4378 4380 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.83893e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.16e-14 panw9=1.2e-14 panw10=0 $X=20140 $Y=59460 $D=111
M9852 4392 4381 4382 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=1.41857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.16e-14 panw9=1.2e-14 panw10=0 $X=20870 $Y=59460 $D=111
M9853 VDD 4385 4392 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30238e-13 as=2.94e-14 pd=8.27387e-07 ps=4.9e-07 nrd=1.6612 nrs=0.375 sa=1.72321e-06 sb=1.08857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=21200 $Y=59460 $D=111
M9854 4385 32 VDD VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.84e-14 as=1.76751e-13 pd=7.4e-07 ps=1.12288e-06 nrd=0.473684 nrs=1.22404 sa=1.18763e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=2.64e-14 panw10=0 $X=21930 $Y=59570 $D=111
M9855 VDD 4382 4385 VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50686e-13 as=6.84e-14 pd=1.39215e-06 ps=7.4e-07 nrd=1.04353 nrs=0.473684 sa=1.45289e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=2.64e-14 panw10=0 $X=22410 $Y=59570 $D=111
M9856 4383 4385 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.18963e-13 pd=1.24e-06 ps=1.09907e-06 nrd=1.06667 nrs=1.32181 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=22850 $Y=60050 $D=111
M9857 VDD 4383 4384 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=23790 $Y=59190 $D=111
M9858 109 4385 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=24270 $Y=59190 $D=111
M9859 4404 801 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=16860 $Y=37880 $D=111
M9860 4396 4398 4404 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=17180 $Y=37880 $D=111
M9861 VDD 68 4396 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=17660 $Y=37880 $D=111
M9862 VDD clk 4395 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=18180 $Y=38470 $D=111
M9863 4398 4395 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=18690 $Y=38610 $D=111
M9864 4406 4395 4396 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=19250 $Y=38110 $D=111
M9865 VDD 4397 4406 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=19570 $Y=38110 $D=111
M9866 4397 4396 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=20110 $Y=38110 $D=111
M9867 4399 4395 4397 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.83893e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.16e-14 panw9=1.2e-14 panw10=0 $X=20940 $Y=37860 $D=111
M9868 4409 4398 4399 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=1.41857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.16e-14 panw9=1.2e-14 panw10=0 $X=21670 $Y=37860 $D=111
M9869 VDD 4402 4409 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30238e-13 as=2.94e-14 pd=8.27387e-07 ps=4.9e-07 nrd=1.6612 nrs=0.375 sa=1.72321e-06 sb=1.08857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=22000 $Y=37860 $D=111
M9870 4402 68 VDD VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.84e-14 as=1.76751e-13 pd=7.4e-07 ps=1.12288e-06 nrd=0.473684 nrs=1.22404 sa=1.18763e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=2.64e-14 panw10=0 $X=22730 $Y=37970 $D=111
M9871 VDD 4399 4402 VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50686e-13 as=6.84e-14 pd=1.39215e-06 ps=7.4e-07 nrd=1.04353 nrs=0.473684 sa=1.45289e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=2.64e-14 panw10=0 $X=23210 $Y=37970 $D=111
M9872 4400 4402 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.18963e-13 pd=1.24e-06 ps=1.09907e-06 nrd=1.06667 nrs=1.32181 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=23650 $Y=38450 $D=111
M9873 VDD 4400 4401 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=24590 $Y=37590 $D=111
M9874 159 4402 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=25070 $Y=37590 $D=111
M9875 4421 226 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=54460 $Y=14640 $D=111
M9876 4413 4415 4421 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=54780 $Y=14640 $D=111
M9877 VDD 202 4413 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=55260 $Y=14640 $D=111
M9878 VDD clk 4412 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=55780 $Y=13910 $D=111
M9879 4415 4412 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=56290 $Y=13910 $D=111
M9880 4423 4412 4413 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=56850 $Y=14410 $D=111
M9881 VDD 4414 4423 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=57170 $Y=14410 $D=111
M9882 4414 4413 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=57710 $Y=14410 $D=111
M9883 4416 4412 4414 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.83893e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.16e-14 panw9=1.2e-14 panw10=0 $X=58540 $Y=14660 $D=111
M9884 4426 4415 4416 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=1.41857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.16e-14 panw9=1.2e-14 panw10=0 $X=59270 $Y=14660 $D=111
M9885 VDD 4419 4426 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30238e-13 as=2.94e-14 pd=8.27387e-07 ps=4.9e-07 nrd=1.6612 nrs=0.375 sa=1.72321e-06 sb=1.08857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=59600 $Y=14660 $D=111
M9886 4419 202 VDD VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.84e-14 as=1.76751e-13 pd=7.4e-07 ps=1.12288e-06 nrd=0.473684 nrs=1.22404 sa=1.18763e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=2.64e-14 panw10=0 $X=60330 $Y=14450 $D=111
M9887 VDD 4416 4419 VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50686e-13 as=6.84e-14 pd=1.39215e-06 ps=7.4e-07 nrd=1.04353 nrs=0.473684 sa=1.45289e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=2.64e-14 panw10=0 $X=60810 $Y=14450 $D=111
M9888 4417 4419 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.18963e-13 pd=1.24e-06 ps=1.09907e-06 nrd=1.06667 nrs=1.32181 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=61250 $Y=14050 $D=111
M9889 VDD 4417 4418 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=62190 $Y=13930 $D=111
M9890 143 4419 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=62670 $Y=13930 $D=111
M9891 4438 261 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=62860 $Y=16280 $D=111
M9892 4430 4432 4438 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=63180 $Y=16280 $D=111
M9893 VDD 299 4430 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=63660 $Y=16280 $D=111
M9894 VDD clk 4429 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=64180 $Y=16870 $D=111
M9895 4432 4429 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=64690 $Y=17010 $D=111
M9896 4440 4429 4430 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=65250 $Y=16510 $D=111
M9897 VDD 4431 4440 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=65570 $Y=16510 $D=111
M9898 4431 4430 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=66110 $Y=16510 $D=111
M9899 4433 4429 4431 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.83893e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.16e-14 panw9=1.2e-14 panw10=0 $X=66940 $Y=16260 $D=111
M9900 4443 4432 4433 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=1.41857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.16e-14 panw9=1.2e-14 panw10=0 $X=67670 $Y=16260 $D=111
M9901 VDD 4436 4443 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30238e-13 as=2.94e-14 pd=8.27387e-07 ps=4.9e-07 nrd=1.6612 nrs=0.375 sa=1.72321e-06 sb=1.08857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=68000 $Y=16260 $D=111
M9902 4436 299 VDD VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.84e-14 as=1.76751e-13 pd=7.4e-07 ps=1.12288e-06 nrd=0.473684 nrs=1.22404 sa=1.18763e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=2.64e-14 panw10=0 $X=68730 $Y=16370 $D=111
M9903 VDD 4433 4436 VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50686e-13 as=6.84e-14 pd=1.39215e-06 ps=7.4e-07 nrd=1.04353 nrs=0.473684 sa=1.45289e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=2.64e-14 panw10=0 $X=69210 $Y=16370 $D=111
M9904 4434 4436 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.18963e-13 pd=1.24e-06 ps=1.09907e-06 nrd=1.06667 nrs=1.32181 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=69650 $Y=16850 $D=111
M9905 VDD 4434 4435 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=70590 $Y=15990 $D=111
M9906 264 4436 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=71070 $Y=15990 $D=111
M9907 4455 827 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=1.302e-13 pd=4.8e-07 ps=1.21e-06 nrd=0.357143 nrs=1.66071 sa=3.7e-07 sb=1.63e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=77260 $Y=23480 $D=111
M9908 4447 4449 4455 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.04e-14 as=2.8e-14 pd=6.4e-07 ps=4.8e-07 nrd=0.642857 nrs=0.357143 sa=6.9e-07 sb=1.31e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=77580 $Y=23480 $D=111
M9909 VDD 303 4447 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.36244e-13 as=5.04e-14 pd=1.13778e-06 ps=6.4e-07 nrd=1.73781 nrs=0.642857 sa=1.17e-06 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=78060 $Y=23480 $D=111
M9910 VDD clk 4446 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.04367e-13 as=1.344e-13 pd=1.70667e-06 ps=1.48e-06 nrd=1.15854 nrs=0.761905 sa=3.2e-07 sb=6.83333e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.44e-14 panw8=0 panw9=0 panw10=0 $X=78580 $Y=24070 $D=111
M9911 4449 4446 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.008e-13 as=1.36244e-13 pd=1.28e-06 ps=1.13778e-06 nrd=1.28571 nrs=1.73781 sa=8.3e-07 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=9.6e-15 panw7=0 panw8=0 panw9=0 panw10=0 $X=79090 $Y=24210 $D=111
M9912 4457 4446 4447 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.8e-14 as=2.1e-13 pd=4.8e-07 ps=2.06e-06 nrd=0.357143 nrs=2.67857 sa=3.6e-07 sb=1.51786e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=79650 $Y=23710 $D=111
M9913 VDD 4448 4457 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.88e-14 as=2.8e-14 pd=7e-07 ps=4.8e-07 nrd=0.75 nrs=0.357143 sa=6.8e-07 sb=1.23214e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=79970 $Y=23710 $D=111
M9914 4448 4447 VDD VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.7945e-13 as=5.88e-14 pd=1.31e-06 ps=7e-07 nrd=2.2889 nrs=0.75 sa=1.22e-06 sb=7.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.4e-14 panw9=9.6e-15 panw10=0 $X=80510 $Y=23710 $D=111
M9915 4450 4446 4448 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.665e-14 as=1.7945e-13 pd=9.4e-07 ps=1.31e-06 nrd=1.23278 nrs=2.2889 sa=7.76786e-07 sb=1.83893e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.16e-14 panw9=1.2e-14 panw10=0 $X=81340 $Y=23460 $D=111
M9916 4460 4449 4450 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.94e-14 as=9.665e-14 pd=4.9e-07 ps=9.4e-07 nrd=0.375 nrs=1.23278 sa=1.42857e-06 sb=1.41857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=2.16e-14 panw9=1.2e-14 panw10=0 $X=82070 $Y=23460 $D=111
M9917 VDD 4453 4460 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.30238e-13 as=2.94e-14 pd=8.27387e-07 ps=4.9e-07 nrd=1.6612 nrs=0.375 sa=1.72321e-06 sb=1.08857e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=3.36e-14 panw10=0 $X=82400 $Y=23460 $D=111
M9918 4453 303 VDD VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.84e-14 as=1.76751e-13 pd=7.4e-07 ps=1.12288e-06 nrd=0.473684 nrs=1.22404 sa=1.18763e-06 sb=7.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=2.64e-14 panw10=0 $X=83130 $Y=23570 $D=111
M9919 VDD 4450 4453 VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.50686e-13 as=6.84e-14 pd=1.39215e-06 ps=7.4e-07 nrd=1.04353 nrs=0.473684 sa=1.45289e-06 sb=2.4e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=1.92e-14 panw9=2.64e-14 panw10=0 $X=83610 $Y=23570 $D=111
M9920 4451 4453 VDD VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=9.6e-14 as=1.18963e-13 pd=1.24e-06 ps=1.09907e-06 nrd=1.06667 nrs=1.32181 sa=2.4e-07 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=1.2e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.68e-14 panw8=0 panw9=0 panw10=0 $X=84050 $Y=24050 $D=111
M9921 VDD 4451 4452 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=8e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=84990 $Y=23190 $D=111
M9922 298 4453 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=8e-07 sb=3.2e-07 sd=0 panw1=0 panw2=3.6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=85470 $Y=23190 $D=111
M9923 4463 22 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.961e-13 as=3.922e-13 pd=1.43e-06 ps=2.86e-06 nrd=0.174528 nrs=0.349057 sa=3.7e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=12580 $Y=30630 $D=111
M9924 VDD 42 4463 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.41646e-13 as=1.961e-13 pd=1.76667e-06 ps=1.43e-06 nrd=0.304064 nrs=0.174528 sa=8.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=13070 $Y=30630 $D=111
M9925 800 4463 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.12554e-13 pd=1.64e-06 ps=2.13333e-06 nrd=0.140625 nrs=0.251803 sa=1.40078e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=13860 $Y=30410 $D=111
M9926 VDD 62 800 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.77313e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=14340 $Y=30410 $D=111
M9927 800 62 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.85563e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=14820 $Y=30410 $D=111
M9928 VDD 4463 800 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=1.93813e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=15300 $Y=30410 $D=111
M9929 4468 215 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.961e-13 as=3.922e-13 pd=1.43e-06 ps=2.86e-06 nrd=0.174528 nrs=0.349057 sa=3.7e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=58980 $Y=64310 $D=111
M9930 VDD 222 4468 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.41646e-13 as=1.961e-13 pd=1.76667e-06 ps=1.43e-06 nrd=0.304064 nrs=0.174528 sa=8.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=59470 $Y=64310 $D=111
M9931 225 4468 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.12554e-13 pd=1.64e-06 ps=2.13333e-06 nrd=0.140625 nrs=0.251803 sa=1.40078e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=60260 $Y=64310 $D=111
M9932 VDD 233 225 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.77313e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=60740 $Y=64310 $D=111
M9933 225 233 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.85563e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=61220 $Y=64310 $D=111
M9934 VDD 4468 225 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=1.93813e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=61700 $Y=64310 $D=111
M9935 4473 265 VDD VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.961e-13 as=3.922e-13 pd=1.43e-06 ps=2.86e-06 nrd=0.174528 nrs=0.349057 sa=3.7e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=71780 $Y=42710 $D=111
M9936 VDD 270 4473 VDD lppfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.41646e-13 as=1.961e-13 pd=1.76667e-06 ps=1.43e-06 nrd=0.304064 nrs=0.174528 sa=8.6e-07 sb=2e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.32e-14 panw10=0 $X=72270 $Y=42710 $D=111
M9937 824 4473 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.12554e-13 pd=1.64e-06 ps=2.13333e-06 nrd=0.140625 nrs=0.251803 sa=1.40078e-06 sb=1.76e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=73060 $Y=42710 $D=111
M9938 VDD 292 824 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.77313e-06 sb=1.28e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=73540 $Y=42710 $D=111
M9939 824 292 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=2.304e-13 pd=1.64e-06 ps=1.64e-06 nrd=0.140625 nrs=0.140625 sa=1.85563e-06 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=74020 $Y=42710 $D=111
M9940 VDD 4473 824 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=2.304e-13 pd=3.2e-06 ps=1.64e-06 nrd=0.25 nrs=0.140625 sa=1.93813e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=74500 $Y=42710 $D=111
M9941 VDD 45 4478 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12667e-13 as=9.6e-14 pd=8.77778e-07 ps=1.24e-06 nrd=1.25185 nrs=1.06667 sa=3.2e-07 sb=1.456e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=12850 $Y=57200 $D=111
M9942 4480 31 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.92933e-13 pd=1.14e-06 ps=2.28222e-06 nrd=0.230769 nrs=0.481481 sa=5.6e-07 sb=1.57692e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=13410 $Y=57200 $D=111
M9943 25 4478 4480 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62584e-13 as=1.404e-13 pd=1.37766e-06 ps=1.14e-06 nrd=0.267233 nrs=0.230769 sa=1.04e-06 sb=1.09692e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=13890 $Y=57200 $D=111
M9944 4479 45 25 VDD lppfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.052e-13 as=1.58416e-13 pd=1.3e-06 ps=1.34234e-06 nrd=0.355263 nrs=0.274265 sa=1.05711e-06 sb=9.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.68e-14 panw10=0 $X=14370 $Y=57440 $D=111
M9945 VDD 4480 4479 VDD lppfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.432e-13 as=2.052e-13 pd=2.16e-06 ps=1.3e-06 nrd=0.421053 nrs=0.355263 sa=1.67763e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.68e-14 panw10=0 $X=15030 $Y=57440 $D=111
M9946 VDD 192 4481 VDD lppfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.12667e-13 as=9.6e-14 pd=8.77778e-07 ps=1.24e-06 nrd=1.25185 nrs=1.06667 sa=3.2e-07 sb=1.456e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=1.08e-14 panw8=0 panw9=0 panw10=0 $X=67250 $Y=35600 $D=111
M9947 4483 231 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.404e-13 as=2.92933e-13 pd=1.14e-06 ps=2.28222e-06 nrd=0.230769 nrs=0.481481 sa=5.6e-07 sb=1.57692e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=67810 $Y=35600 $D=111
M9948 820 4481 4483 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.62584e-13 as=1.404e-13 pd=1.37766e-06 ps=1.14e-06 nrd=0.267233 nrs=0.230769 sa=1.04e-06 sb=1.09692e-06 sd=0 panw1=0 panw2=0 panw3=1.2e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=2.04e-14 panw10=0 $X=68290 $Y=35600 $D=111
M9949 4482 192 820 VDD lppfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.052e-13 as=1.58416e-13 pd=1.3e-06 ps=1.34234e-06 nrd=0.355263 nrs=0.274265 sa=1.05711e-06 sb=9.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.68e-14 panw10=0 $X=68770 $Y=35840 $D=111
M9950 VDD 4483 4482 VDD lppfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.432e-13 as=2.052e-13 pd=2.16e-06 ps=1.3e-06 nrd=0.421053 nrs=0.355263 sa=1.67763e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.04e-14 panw8=2.4e-14 panw9=4.68e-14 panw10=0 $X=69430 $Y=35840 $D=111
M9951 VDD 60 4484 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.57647e-14 as=1.008e-13 pd=7.57647e-07 ps=1.28e-06 nrd=0.966387 nrs=1.28571 sa=3.6e-07 sb=1.25714e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=9.6e-15 panw9=0 panw10=0 $X=14960 $Y=67110 $D=111
M9952 4486 54 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16615e-13 as=1.08235e-13 pd=1.12821e-06 ps=1.08235e-06 nrd=0.728846 nrs=0.676471 sa=7.96e-07 sb=5.66e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=15600 $Y=66990 $D=111
M9953 41 4484 4486 VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22477e-13 as=1.10785e-13 pd=1.10103e-06 ps=1.07179e-06 nrd=0.848178 nrs=0.767206 sa=5.64737e-07 sb=4.93158e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=9.6e-15 panw8=0 panw9=0 panw10=0 $X=16120 $Y=67310 $D=111
M9954 4485 60 41 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=1.28923e-13 pd=1.31e-06 ps=1.15897e-06 nrd=1.1375 nrs=0.805769 sa=6.8e-07 sb=4.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=16670 $Y=66990 $D=111
M9955 4485 4486 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=6.4e-14 pd=1.31e-06 ps=7.2e-07 nrd=1.1375 nrs=0.4 sa=5.2e-07 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=4.8e-14 $X=16870 $Y=66440 $D=111
M9956 VDD 116 4487 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.57647e-14 as=1.008e-13 pd=7.57647e-07 ps=1.28e-06 nrd=0.966387 nrs=1.28571 sa=3.6e-07 sb=1.25714e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=9.6e-15 panw9=0 panw10=0 $X=34160 $Y=16710 $D=111
M9957 4489 118 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16615e-13 as=1.08235e-13 pd=1.12821e-06 ps=1.08235e-06 nrd=0.728846 nrs=0.676471 sa=7.96e-07 sb=5.66e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=34800 $Y=16590 $D=111
M9958 122 4487 4489 VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22477e-13 as=1.10785e-13 pd=1.10103e-06 ps=1.07179e-06 nrd=0.848178 nrs=0.767206 sa=5.64737e-07 sb=4.93158e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=9.6e-15 panw8=0 panw9=0 panw10=0 $X=35320 $Y=16910 $D=111
M9959 4488 116 122 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=1.28923e-13 pd=1.31e-06 ps=1.15897e-06 nrd=1.1375 nrs=0.805769 sa=6.8e-07 sb=4.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=35870 $Y=16590 $D=111
M9960 4488 4489 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=6.4e-14 pd=1.31e-06 ps=7.2e-07 nrd=1.1375 nrs=0.4 sa=6.955e-07 sb=8.3e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=4.8e-14 $X=36070 $Y=16040 $D=111
M9961 VDD 259 4490 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.57647e-14 as=1.008e-13 pd=7.57647e-07 ps=1.28e-06 nrd=0.966387 nrs=1.28571 sa=3.6e-07 sb=1.25714e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=9.6e-15 panw9=0 panw10=0 $X=66560 $Y=21410 $D=111
M9962 4492 281 VDD VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.16615e-13 as=1.08235e-13 pd=1.12821e-06 ps=1.08235e-06 nrd=0.728846 nrs=0.676471 sa=7.96e-07 sb=5.66e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=67200 $Y=21410 $D=111
M9963 257 4490 4492 VDD lppfet w=3.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.22477e-13 as=1.10785e-13 pd=1.10103e-06 ps=1.07179e-06 nrd=0.848178 nrs=0.767206 sa=5.64737e-07 sb=4.93158e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=9.6e-15 panw8=0 panw9=0 panw10=0 $X=67720 $Y=21110 $D=111
M9964 4491 259 257 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.82e-13 as=1.28923e-13 pd=1.31e-06 ps=1.15897e-06 nrd=1.1375 nrs=0.805769 sa=6.8e-07 sb=4.8e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=2.4e-14 panw8=2.4e-14 panw9=0 panw10=0 $X=68270 $Y=21410 $D=111
M9965 VDD 4492 4491 VDD lppfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.4e-14 as=1.82e-13 pd=7.2e-07 ps=1.31e-06 nrd=0.4 nrs=1.1375 sa=8.3e-07 sb=1.556e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=4.8e-14 $X=68470 $Y=22240 $D=111
M9966 VDD 39 4493 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.11724e-13 as=3.712e-13 pd=1.54017e-06 ps=2.96e-06 nrd=0.157346 nrs=0.275862 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=16260 $Y=16050 $D=111
M9967 29 46 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.196e-13 as=2.22676e-13 pd=1.58e-06 ps=1.61983e-06 nrd=0.147541 nrs=0.149607 sa=7.74426e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=16740 $Y=15990 $D=111
M9968 VDD 4493 29 VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.196e-13 as=2.196e-13 pd=1.58e-06 ps=1.58e-06 nrd=0.147541 nrs=0.147541 sa=1.25443e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=17220 $Y=15990 $D=111
M9969 29 4493 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.196e-13 as=2.196e-13 pd=1.58e-06 ps=1.58e-06 nrd=0.147541 nrs=0.147541 sa=1.73443e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=17700 $Y=15990 $D=111
M9970 VDD 46 29 VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.196e-13 pd=3.08e-06 ps=1.58e-06 nrd=0.262295 nrs=0.147541 sa=1.98623e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=18180 $Y=15990 $D=111
M9971 VDD 162 4497 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.11724e-13 as=3.712e-13 pd=1.54017e-06 ps=2.96e-06 nrd=0.157346 nrs=0.275862 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=53460 $Y=42790 $D=111
M9972 206 135 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.196e-13 as=2.22676e-13 pd=1.58e-06 ps=1.61983e-06 nrd=0.147541 nrs=0.149607 sa=7.74426e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=53940 $Y=42790 $D=111
M9973 VDD 4497 206 VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.196e-13 as=2.196e-13 pd=1.58e-06 ps=1.58e-06 nrd=0.147541 nrs=0.147541 sa=1.25443e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=54420 $Y=42790 $D=111
M9974 206 4497 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.196e-13 as=2.196e-13 pd=1.58e-06 ps=1.58e-06 nrd=0.147541 nrs=0.147541 sa=1.73443e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=54900 $Y=42790 $D=111
M9975 VDD 135 206 VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.196e-13 pd=3.08e-06 ps=1.58e-06 nrd=0.262295 nrs=0.147541 sa=1.98623e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=55380 $Y=42790 $D=111
M9976 VDD 205 4501 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.11724e-13 as=3.712e-13 pd=1.54017e-06 ps=2.96e-06 nrd=0.157346 nrs=0.275862 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=54660 $Y=23250 $D=111
M9977 207 204 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.196e-13 as=2.22676e-13 pd=1.58e-06 ps=1.61983e-06 nrd=0.147541 nrs=0.149607 sa=7.74426e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=55140 $Y=23190 $D=111
M9978 VDD 4501 207 VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.196e-13 as=2.196e-13 pd=1.58e-06 ps=1.58e-06 nrd=0.147541 nrs=0.147541 sa=1.25443e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=55620 $Y=23190 $D=111
M9979 207 4501 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.196e-13 as=2.196e-13 pd=1.58e-06 ps=1.58e-06 nrd=0.147541 nrs=0.147541 sa=1.73443e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=56100 $Y=23190 $D=111
M9980 VDD 204 207 VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.196e-13 pd=3.08e-06 ps=1.58e-06 nrd=0.262295 nrs=0.147541 sa=1.98623e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=56580 $Y=23190 $D=111
M9981 VDD 135 4505 VDD lppfet w=1.16e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.11724e-13 as=3.712e-13 pd=1.54017e-06 ps=2.96e-06 nrd=0.157346 nrs=0.275862 sa=3.2e-07 sb=2e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.68e-14 $X=61460 $Y=42790 $D=111
M9982 216 162 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.196e-13 as=2.22676e-13 pd=1.58e-06 ps=1.61983e-06 nrd=0.147541 nrs=0.149607 sa=7.74426e-07 sb=1.76e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=61940 $Y=42790 $D=111
M9983 VDD 4505 216 VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.196e-13 as=2.196e-13 pd=1.58e-06 ps=1.58e-06 nrd=0.147541 nrs=0.147541 sa=1.25443e-06 sb=1.28e-06 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=62420 $Y=42790 $D=111
M9984 216 4505 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.196e-13 as=2.196e-13 pd=1.58e-06 ps=1.58e-06 nrd=0.147541 nrs=0.147541 sa=1.73443e-06 sb=8e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=62900 $Y=42790 $D=111
M9985 VDD 162 216 VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.904e-13 as=2.196e-13 pd=3.08e-06 ps=1.58e-06 nrd=0.262295 nrs=0.147541 sa=1.98623e-06 sb=3.2e-07 sd=0 panw1=0 panw2=0 panw3=2.4e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=63380 $Y=42790 $D=111
M9986 4510 4511 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.11812e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=20020 $Y=21110 $D=111
M9987 VDD 4511 4510 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.348e-13 as=2.304e-13 pd=2.03e-06 ps=1.64e-06 nrd=0.143311 nrs=0.140625 sa=8e-07 sb=6.38125e-07 sd=0 panw1=0 panw2=4.5e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.31e-14 $X=20500 $Y=21110 $D=111
M9988 4509 106 VDD VDD lppfet w=1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.2e-13 as=1.83437e-13 pd=2.64e-06 ps=1.58594e-06 nrd=0.32 nrs=0.183437 sa=1.2192e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.72e-14 panw10=0 $X=20940 $Y=21090 $D=111
M9989 4510 106 126 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=4.064e-13 pd=1.63e-06 ps=3.18e-06 nrd=0.141732 nrs=0.251969 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=21960 $Y=21140 $D=111
M9990 126 106 4510 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.54e-13 as=2.286e-13 pd=1.67e-06 ps=1.63e-06 nrd=0.15748 nrs=0.141732 sa=8e-07 sb=1.44e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=22440 $Y=21140 $D=111
M9991 4511 4509 126 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.54e-13 pd=1.63e-06 ps=1.67e-06 nrd=0.141732 nrs=0.15748 sa=1.32e-06 sb=9.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=22960 $Y=21140 $D=111
M9992 126 4509 4511 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.588e-13 as=2.286e-13 pd=3.42e-06 ps=1.63e-06 nrd=0.346457 nrs=0.141732 sa=1.8e-06 sb=4.4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=23440 $Y=21140 $D=111
M9993 4512 106 VDD VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.05e-13 as=1.56243e-13 pd=9.2e-07 ps=1.05291e-06 nrd=0.42 nrs=0.624974 sa=2.4e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=24540 $Y=21140 $D=111
M9994 VDD 100 4512 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.56243e-13 as=1.05e-13 pd=1.05291e-06 ps=9.2e-07 nrd=0.624974 nrs=0.42 sa=7.8e-07 sb=1.72e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=25080 $Y=21140 $D=111
M9995 4511 100 VDD VDD lppfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.16e-13 as=3.74984e-13 pd=1.56e-06 ps=2.52698e-06 nrd=0.15 nrs=0.260406 sa=9.42333e-07 sb=1.28e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.56e-14 $X=25520 $Y=21140 $D=111
M9996 VDD 100 4511 VDD lppfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.16e-13 as=2.16e-13 pd=1.56e-06 ps=1.56e-06 nrd=0.15 nrs=0.15 sa=1.42233e-06 sb=8e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.56e-14 $X=26000 $Y=21140 $D=111
M9997 4511 100 VDD VDD lppfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.84e-13 as=2.16e-13 pd=3.04e-06 ps=1.56e-06 nrd=0.266667 nrs=0.15 sa=1.77333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.56e-14 $X=26480 $Y=21140 $D=111
M9998 90 4512 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.096e-13 pd=3.2e-06 ps=3.2e-06 nrd=0.25 nrs=0.25 sa=3.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=27470 $Y=21110 $D=111
M9999 4515 4516 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.304e-13 as=4.096e-13 pd=1.64e-06 ps=3.2e-06 nrd=0.140625 nrs=0.25 sa=3.2e-07 sb=1.11812e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=52420 $Y=35510 $D=111
M10000 VDD 4516 4515 VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.348e-13 as=2.304e-13 pd=2.03e-06 ps=1.64e-06 nrd=0.143311 nrs=0.140625 sa=8e-07 sb=6.38125e-07 sd=0 panw1=0 panw2=4.5e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.31e-14 $X=52900 $Y=35510 $D=111
M10001 4514 224 VDD VDD lppfet w=1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.2e-13 as=1.83437e-13 pd=2.64e-06 ps=1.58594e-06 nrd=0.32 nrs=0.183437 sa=1.2192e-06 sb=3.2e-07 sd=0 panw1=0 panw2=4.8e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=3.72e-14 panw10=0 $X=53340 $Y=35490 $D=111
M10002 4515 224 150 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=4.064e-13 pd=1.63e-06 ps=3.18e-06 nrd=0.141732 nrs=0.251969 sa=3.2e-07 sb=1.92e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=54360 $Y=35540 $D=111
M10003 150 224 4515 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.54e-13 as=2.286e-13 pd=1.67e-06 ps=1.63e-06 nrd=0.15748 nrs=0.141732 sa=8e-07 sb=1.44e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=54840 $Y=35540 $D=111
M10004 4516 4514 150 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=2.54e-13 pd=1.63e-06 ps=1.67e-06 nrd=0.141732 nrs=0.15748 sa=1.32e-06 sb=9.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=55360 $Y=35540 $D=111
M10005 150 4514 4516 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=5.588e-13 as=2.286e-13 pd=3.42e-06 ps=1.63e-06 nrd=0.346457 nrs=0.141732 sa=1.8e-06 sb=4.4e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.4e-14 $X=55840 $Y=35540 $D=111
M10006 4517 224 VDD VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.05e-13 as=1.56243e-13 pd=9.2e-07 ps=1.05291e-06 nrd=0.42 nrs=0.624974 sa=2.4e-07 sb=2e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=56940 $Y=35540 $D=111
M10007 VDD 159 4517 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.56243e-13 as=1.05e-13 pd=1.05291e-06 ps=9.2e-07 nrd=0.624974 nrs=0.42 sa=7.8e-07 sb=1.72e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=3.6e-15 panw9=0 panw10=0 $X=57480 $Y=35540 $D=111
M10008 4516 159 VDD VDD lppfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.16e-13 as=3.74984e-13 pd=1.56e-06 ps=2.52698e-06 nrd=0.15 nrs=0.260406 sa=9.42333e-07 sb=1.28e-06 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.56e-14 $X=57920 $Y=35540 $D=111
M10009 VDD 159 4516 VDD lppfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.16e-13 as=2.16e-13 pd=1.56e-06 ps=1.56e-06 nrd=0.15 nrs=0.15 sa=1.42233e-06 sb=8e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.56e-14 $X=58400 $Y=35540 $D=111
M10010 4516 159 VDD VDD lppfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=3.84e-13 as=2.16e-13 pd=3.04e-06 ps=1.56e-06 nrd=0.266667 nrs=0.15 sa=1.77333e-06 sb=3.2e-07 sd=0 panw1=0 panw2=2.4e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.56e-14 $X=58880 $Y=35540 $D=111
M10011 223 4517 VDD VDD lppfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.096e-13 as=4.096e-13 pd=3.2e-06 ps=3.2e-06 nrd=0.25 nrs=0.25 sa=3.2e-07 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.16e-14 $X=59870 $Y=35510 $D=111
M10012 VDD 101 4519 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.272e-14 as=9.24e-14 pd=6.56e-07 ps=1.22e-06 nrd=0.8 nrs=1.17857 sa=3.3e-07 sb=1.37e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=1.56e-14 panw9=0 panw10=0 $X=32020 $Y=31060 $D=111
M10013 102 78 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.56e-14 as=9.408e-14 pd=7.8e-07 ps=9.84e-07 nrd=0.428571 nrs=0.533333 sa=6.73333e-07 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=32540 $Y=30920 $D=111
M10014 VDD 4519 102 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.453e-13 as=7.56e-14 pd=2.2e-06 ps=7.8e-07 nrd=1.39059 nrs=0.428571 sa=1.15333e-06 sb=3.7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=33020 $Y=30920 $D=111
M10015 VDD 217 4521 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=6.272e-14 as=9.24e-14 pd=6.56e-07 ps=1.22e-06 nrd=0.8 nrs=1.17857 sa=3.3e-07 sb=1.37e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=1.56e-14 panw9=0 panw10=0 $X=52420 $Y=23860 $D=111
M10016 814 113 VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=7.56e-14 as=9.408e-14 pd=7.8e-07 ps=9.84e-07 nrd=0.428571 nrs=0.533333 sa=6.73333e-07 sb=8.5e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=52940 $Y=23720 $D=111
M10017 VDD 4521 814 VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.453e-13 as=7.56e-14 pd=2.2e-06 ps=7.8e-07 nrd=1.39059 nrs=0.428571 sa=1.15333e-06 sb=3.7e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=1.8e-14 panw8=2.4e-14 panw9=8.4e-15 panw10=0 $X=53420 $Y=23720 $D=111
M10018 VDD data_in[0] 4523 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.06026e-13 as=2.56e-13 pd=1.36851e-06 ps=2.24e-06 nrd=0.321915 nrs=0.4 sa=3.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.2e-13 panw9=1.2e-14 panw10=0 $X=8910 $Y=16490 $D=111
M10019 101 4523 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=3.27066e-13 pd=1.63e-06 ps=2.17251e-06 nrd=0.141732 nrs=0.202781 sa=6.87559e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.728e-13 $X=9470 $Y=16020 $D=111
M10020 VDD 4523 101 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.43435e-13 as=2.286e-13 pd=3.16271e-06 ps=1.63e-06 nrd=0.27493 nrs=0.141732 sa=1.16756e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=1.601e-13 $X=9950 $Y=16020 $D=111
M10021 VDD weight_in[6] 4524 VDD lppfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.06026e-13 as=2.56e-13 pd=1.36851e-06 ps=2.24e-06 nrd=0.321915 nrs=0.4 sa=3.2e-07 sb=1.4e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=1.2e-14 panw10=0 $X=46510 $Y=74090 $D=111
M10022 195 4524 VDD VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.286e-13 as=3.27066e-13 pd=1.63e-06 ps=2.17251e-06 nrd=0.141732 nrs=0.202781 sa=6.87559e-07 sb=8.4e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.04e-14 $X=47070 $Y=73620 $D=111
M10023 VDD 4524 195 VDD lppfet w=1.27e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=4.43435e-13 as=2.286e-13 pd=3.16271e-06 ps=1.63e-06 nrd=0.27493 nrs=0.141732 sa=1.16756e-06 sb=3.6e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=2.4e-14 panw9=4.8e-14 panw10=2.04e-14 $X=47550 $Y=73620 $D=111
M10024 VDD data_in[7] 4525 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07368e-13 as=1.6e-13 pd=9.12281e-07 ps=1.64e-06 nrd=0.429474 nrs=0.64 sa=3.2e-07 sb=1.32e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=10840 $Y=57110 $D=111
M10025 186 4525 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.37432e-13 pd=1e-06 ps=1.16772e-06 nrd=0.28125 nrs=0.335526 sa=7.2625e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=11360 $Y=57110 $D=111
M10026 VDD 4525 186 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.152e-13 pd=1.92e-06 ps=1e-06 nrd=0.5 nrs=0.28125 sa=1.20625e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=11840 $Y=57110 $D=111
M10027 VDD weight_in[3] 4526 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.07368e-13 as=1.6e-13 pd=9.12281e-07 ps=1.64e-06 nrd=0.429474 nrs=0.64 sa=3.2e-07 sb=1.32e-06 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=0 panw9=0 panw10=0 $X=34440 $Y=64310 $D=111
M10028 111 4526 VDD VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=1.152e-13 as=1.37432e-13 pd=1e-06 ps=1.16772e-06 nrd=0.28125 nrs=0.335526 sa=7.2625e-07 sb=8e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=34960 $Y=64310 $D=111
M10029 VDD 4526 111 VDD lppfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 ad=2.048e-13 as=1.152e-13 pd=1.92e-06 ps=1e-06 nrd=0.5 nrs=0.28125 sa=1.20625e-06 sb=3.2e-07 sd=0 panw1=0 panw2=6e-15 panw3=6e-15 panw4=6e-15 panw5=6e-15 panw6=1.2e-14 panw7=2.4e-14 panw8=1.68e-14 panw9=0 panw10=0 $X=35440 $Y=64310 $D=111
D10030 VSS VDD diodenwx AREA=7.15473e-10 perim=0.00037152 t3well=0 $X=8060 $Y=71210 $D=474
D10031 VSS VDD diodenwx AREA=7.1777e-10 perim=0.00037048 t3well=0 $X=8060 $Y=28010 $D=474
D10032 VSS VDD diodenwx AREA=7.17032e-10 perim=0.00037146 t3well=0 $X=8060 $Y=13610 $D=474
D10033 VSS VDD diodenwx AREA=7.11911e-10 perim=0.00037268 t3well=0 $X=8060 $Y=64010 $D=474
D10034 VSS VDD diodenwx AREA=7.17389e-10 perim=0.0003708 t3well=0 $X=8060 $Y=20810 $D=474
D10035 VSS VDD diodenwx AREA=7.15089e-10 perim=0.0003717 t3well=0 $X=8060 $Y=42410 $D=474
D10036 VSS VDD diodenwx AREA=7.14297e-10 perim=0.00037244 t3well=0 $X=8060 $Y=35210 $D=474
D10037 VSS VDD diodenwx AREA=7.18004e-10 perim=0.00037086 t3well=0 $X=8060 $Y=56810 $D=474
D10038 VSS VDD diodenwx AREA=7.15227e-10 perim=0.0003717 t3well=0 $X=8060 $Y=49610 $D=474
D10039 VSS VDD diodenwx AREA=4.31825e-10 perim=0.00036614 t3well=0 $X=8060 $Y=8000 $D=474
.ENDS
***************************************
