##
## LEF for PtnCells ;
## created by Innovus v19.10-p002_1 on Sat Apr  9 14:54:28 2022
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO PE
  CLASS BLOCK ;
  SIZE 196.800000 BY 85.200000 ;
  FOREIGN PE 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 11.900000 84.600000 12.100000 85.200000 ;
    END
  END clk
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 16.900000 84.600000 17.100000 85.200000 ;
    END
  END rst_n
  PIN fire_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.900000 84.600000 55.100000 85.200000 ;
    END
  END fire_in
  PIN weight_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 47.400000 84.600000 47.600000 85.200000 ;
    END
  END weight_in[7]
  PIN weight_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 43.900000 84.600000 44.100000 85.200000 ;
    END
  END weight_in[6]
  PIN weight_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 40.400000 84.600000 40.600000 85.200000 ;
    END
  END weight_in[5]
  PIN weight_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 36.900000 84.600000 37.100000 85.200000 ;
    END
  END weight_in[4]
  PIN weight_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 33.400000 84.600000 33.600000 85.200000 ;
    END
  END weight_in[3]
  PIN weight_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 29.900000 84.600000 30.100000 85.200000 ;
    END
  END weight_in[2]
  PIN weight_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 26.400000 84.600000 26.600000 85.200000 ;
    END
  END weight_in[1]
  PIN weight_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 22.900000 84.600000 23.100000 85.200000 ;
    END
  END weight_in[0]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 54.900000 0.600000 55.100000 ;
    END
  END data_in[7]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 49.900000 0.600000 50.100000 ;
    END
  END data_in[6]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 44.900000 0.600000 45.100000 ;
    END
  END data_in[5]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 39.900000 0.600000 40.100000 ;
    END
  END data_in[4]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 34.900000 0.600000 35.100000 ;
    END
  END data_in[3]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 29.900000 0.600000 30.100000 ;
    END
  END data_in[2]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 24.900000 0.600000 25.100000 ;
    END
  END data_in[1]
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 19.900000 0.600000 20.100000 ;
    END
  END data_in[0]
  PIN fire_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.900000 0.000000 55.100000 0.600000 ;
    END
  END fire_out
  PIN weight_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.400000 0.000000 47.600000 0.600000 ;
    END
  END weight_out[7]
  PIN weight_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.900000 0.000000 44.100000 0.600000 ;
    END
  END weight_out[6]
  PIN weight_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.400000 0.000000 40.600000 0.600000 ;
    END
  END weight_out[5]
  PIN weight_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.900000 0.000000 37.100000 0.600000 ;
    END
  END weight_out[4]
  PIN weight_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.400000 0.000000 33.600000 0.600000 ;
    END
  END weight_out[3]
  PIN weight_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.900000 0.000000 30.100000 0.600000 ;
    END
  END weight_out[2]
  PIN weight_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.400000 0.000000 26.600000 0.600000 ;
    END
  END weight_out[1]
  PIN weight_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.900000 0.000000 23.100000 0.600000 ;
    END
  END weight_out[0]
  PIN data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.200000 54.900000 196.800000 55.100000 ;
    END
  END data_out[7]
  PIN data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.200000 49.900000 196.800000 50.100000 ;
    END
  END data_out[6]
  PIN data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.200000 44.900000 196.800000 45.100000 ;
    END
  END data_out[5]
  PIN data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.200000 39.900000 196.800000 40.100000 ;
    END
  END data_out[4]
  PIN data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.200000 34.900000 196.800000 35.100000 ;
    END
  END data_out[3]
  PIN data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.200000 29.900000 196.800000 30.100000 ;
    END
  END data_out[2]
  PIN data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.200000 24.900000 196.800000 25.100000 ;
    END
  END data_out[1]
  PIN data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.200000 19.900000 196.800000 20.100000 ;
    END
  END data_out[0]
  PIN result[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.400000 0.000000 178.600000 0.600000 ;
    END
  END result[31]
  PIN result[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.900000 0.000000 175.100000 0.600000 ;
    END
  END result[30]
  PIN result[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.400000 0.000000 171.600000 0.600000 ;
    END
  END result[29]
  PIN result[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.900000 0.000000 168.100000 0.600000 ;
    END
  END result[28]
  PIN result[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.400000 0.000000 164.600000 0.600000 ;
    END
  END result[27]
  PIN result[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.900000 0.000000 161.100000 0.600000 ;
    END
  END result[26]
  PIN result[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.400000 0.000000 157.600000 0.600000 ;
    END
  END result[25]
  PIN result[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.900000 0.000000 154.100000 0.600000 ;
    END
  END result[24]
  PIN result[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.400000 0.000000 150.600000 0.600000 ;
    END
  END result[23]
  PIN result[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.900000 0.000000 147.100000 0.600000 ;
    END
  END result[22]
  PIN result[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.400000 0.000000 143.600000 0.600000 ;
    END
  END result[21]
  PIN result[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.900000 0.000000 140.100000 0.600000 ;
    END
  END result[20]
  PIN result[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.400000 0.000000 136.600000 0.600000 ;
    END
  END result[19]
  PIN result[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.900000 0.000000 133.100000 0.600000 ;
    END
  END result[18]
  PIN result[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.400000 0.000000 129.600000 0.600000 ;
    END
  END result[17]
  PIN result[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.900000 0.000000 126.100000 0.600000 ;
    END
  END result[16]
  PIN result[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.400000 0.000000 122.600000 0.600000 ;
    END
  END result[15]
  PIN result[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.900000 0.000000 119.100000 0.600000 ;
    END
  END result[14]
  PIN result[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.400000 0.000000 115.600000 0.600000 ;
    END
  END result[13]
  PIN result[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.900000 0.000000 112.100000 0.600000 ;
    END
  END result[12]
  PIN result[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.400000 0.000000 108.600000 0.600000 ;
    END
  END result[11]
  PIN result[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.900000 0.000000 105.100000 0.600000 ;
    END
  END result[10]
  PIN result[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.400000 0.000000 101.600000 0.600000 ;
    END
  END result[9]
  PIN result[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.900000 0.000000 98.100000 0.600000 ;
    END
  END result[8]
  PIN result[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.400000 0.000000 94.600000 0.600000 ;
    END
  END result[7]
  PIN result[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.900000 0.000000 91.100000 0.600000 ;
    END
  END result[6]
  PIN result[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.400000 0.000000 87.600000 0.600000 ;
    END
  END result[5]
  PIN result[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.900000 0.000000 84.100000 0.600000 ;
    END
  END result[4]
  PIN result[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.400000 0.000000 80.600000 0.600000 ;
    END
  END result[3]
  PIN result[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.900000 0.000000 77.100000 0.600000 ;
    END
  END result[2]
  PIN result[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.400000 0.000000 73.600000 0.600000 ;
    END
  END result[1]
  PIN result[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.900000 0.000000 70.100000 0.600000 ;
    END
  END result[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M3 ;
        RECT 1.200000 1.200000 195.600000 3.600000 ;
        RECT 1.200000 81.600000 195.600000 84.000000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M3 ;
        RECT 4.800000 4.800000 192.000000 7.200000 ;
        RECT 4.800000 78.000000 192.000000 80.400000 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 196.800000 85.200000 ;
    LAYER M2 ;
      RECT 0.000000 57.020000 196.800000 85.200000 ;
      RECT 0.000000 52.980000 194.280000 57.020000 ;
      RECT 0.000000 52.020000 196.800000 52.980000 ;
      RECT 0.000000 47.980000 194.280000 52.020000 ;
      RECT 0.000000 47.020000 196.800000 47.980000 ;
      RECT 0.000000 42.980000 194.280000 47.020000 ;
      RECT 0.000000 42.020000 196.800000 42.980000 ;
      RECT 0.000000 37.980000 194.280000 42.020000 ;
      RECT 0.000000 37.020000 196.800000 37.980000 ;
      RECT 0.000000 32.980000 194.280000 37.020000 ;
      RECT 0.000000 32.020000 196.800000 32.980000 ;
      RECT 0.000000 27.980000 194.280000 32.020000 ;
      RECT 0.000000 27.020000 196.800000 27.980000 ;
      RECT 0.000000 22.980000 194.280000 27.020000 ;
      RECT 0.000000 22.020000 196.800000 22.980000 ;
      RECT 0.000000 17.980000 194.280000 22.020000 ;
      RECT 0.000000 2.520000 196.800000 17.980000 ;
      RECT 180.520000 0.000000 196.800000 2.520000 ;
      RECT 57.020000 0.000000 67.980000 2.520000 ;
      RECT 49.520000 0.000000 52.980000 2.520000 ;
      RECT 0.000000 0.000000 20.980000 2.520000 ;
    LAYER M3 ;
      RECT 193.920000 76.080000 196.800000 79.680000 ;
      RECT 0.000000 76.080000 2.880000 79.680000 ;
      RECT 0.000000 57.020000 196.800000 76.080000 ;
      RECT 2.520000 52.980000 196.800000 57.020000 ;
      RECT 0.000000 52.020000 196.800000 52.980000 ;
      RECT 2.520000 47.980000 196.800000 52.020000 ;
      RECT 0.000000 47.020000 196.800000 47.980000 ;
      RECT 2.520000 42.980000 196.800000 47.020000 ;
      RECT 0.000000 42.020000 196.800000 42.980000 ;
      RECT 2.520000 37.980000 196.800000 42.020000 ;
      RECT 0.000000 37.020000 196.800000 37.980000 ;
      RECT 2.520000 32.980000 196.800000 37.020000 ;
      RECT 0.000000 32.020000 196.800000 32.980000 ;
      RECT 2.520000 27.980000 196.800000 32.020000 ;
      RECT 0.000000 27.020000 196.800000 27.980000 ;
      RECT 2.520000 22.980000 196.800000 27.020000 ;
      RECT 0.000000 22.020000 196.800000 22.980000 ;
      RECT 2.520000 17.980000 196.800000 22.020000 ;
      RECT 0.000000 9.120000 196.800000 17.980000 ;
      RECT 193.920000 5.520000 196.800000 9.120000 ;
      RECT 0.000000 5.520000 2.880000 9.120000 ;
  END
END PE

END LIBRARY
